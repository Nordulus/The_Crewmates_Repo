PK   l�WW5O*@?B  �{    cirkitFile.json�}�7��_����J;]m$�zi�!ٚY�ؖ���\��`�S�E��ْ��o?��h�$��A�MXaK�U�ćD"x$~�Xf���X,��jy;[�/Qxy�&[�������f6��������ţ�����כ*ȗUV���T�J�L� &��k$uZ$�:�D�XM�T\<������MAL���KAL%���*6.1�l\
b�1p)�id(�_,��,��|5�eL2+��.r�TA�U@q��"����i|������o�e��f���Oo��r��5�W��͉��I��I�s��e6'a7'e8��Q��#�DL&�lS*��RN|#D��"�t�4��46	�B�d]r��7�r%#��:��R�mQ�u��%��#>	��k��O ��86	���6	��߰I��o$��I�(�M ��9lW���A�םl7ΐ	��J��)�E)��J�NW��%a6@�́�6	��j(�u�=S�)��+��R��Ep[�7q�o��$
��c�0(�&�M ��l?<`�S��$
�=`�0(����A��$
�"�f#C 8_cZ���l_�u�2�⺨�@��]Ui��iT����e�G�Ts��W�l_��I|�SNg*fg�|��&aP�?��A���l_��I|��&aP ��;�kl6	���v�$
��e�0(�j�MBL#��d�0(���M ������p�߮�u]WyRu�$Ƹ����\Y�Q�dEV*���:�$����<��[7��'B�; �GGXt�E'��;��aщ���NayEGXt&���NcyEGXt�s��.�����茏��]��a�leE�.vo�٦�c�m�m�UɰOz�`��w�#��|����;(:¢����94n 0>�;�U�_'v�ⅷn�4�ɮN��b�d�]�V����A��_a��ݪ�8���#0��}��u"�:	���u��dW'b�+�j_p��m����`�����=<�8���#0>{��?p��G`|��xb{a��=j�xU	�����!)0��+K�%p�#�яG?X|�g����~�������ʄ�G`|�0 ��������1F0�����������s�q�[�"p�yLvu��R��G?����Av怣�~���Ϟ���`���^�:�G�(�R��G=�c����إ��W�w�����c/��8���#0>{��?p��G`|��:���������z0������� `���~�����4 ��`���ƀ�G?X|�g�H���~����=���f*/BU �ցN�,HK��C��i"Ҹ�*�^�#'^7��;�W�I7ͦ��t����)������&J�} 
}"
2ip��N�n/8d��;��ɱ�d8��������l:0�����D>`��#.,>�)���G\X|�g3 a��#.,>㳹���G\X|�g�N������������`�Q��P�)y7�M�|Bp���w6��ˮئ��h`֣3I�SI�יBp���,>�����;�Qb�wn�4�i�U��)LX|�g�������Ϧ=��/LX|�g6������Ϧ���%p�N#p��m�^�Hf�S������y;9��U#��D�]�e@i�3�y;��K}y2#N�f�Jpj�^"��9cIp9�Y��zbuD�سnB�T��%��P�~�� �K>�~��">��v��߷3w��$LCֹ�r��LS�\�x���ȓCwq�m0bUr������[q�Z���9U��\�ȑU�����Dq���b^��Tu̪��W:����i�:7���i�T�rк��8X�m�S�9 �"�u�TU�2
��� /T�qT�:�Z�A=�T�qq�yȸ8^t�󯅋{�x�ɰ92�qsĐ�q"F�C�VEy��<	�����E�gF�Fa��,/�H�G��>֢N�+QG��1%�z�ѽ�T=�+8�W���|G��S�����^q���+N�	��!g�ճcT=��zv���cV��L��i�����Z�]ê�q�
�%�4(��Ļ[UP5�YR2j��ڇT�S��!�uIIid>�ei\�BƁ*E���S}��p���������Qɺ�)��tX�AZYjuQ�u(��#��>���0�"�e�GQ���k� �QTB�TuX���N��w�|�.2UGƪ��N]���Z�AH��B�"O��1�χ�;}ހ��|?]-���z��x�g��4��_D���3�A��p�DHX�c�	��1�@��5D B�"!�"jUIX�Q�B[B����h��(����g~�%(D)J�@��5ՆR]SE�6�D�`z�$J���	��Q��E�R�5L{S�'���&O0N �K0J�Y�a�iq��q%�lO 9�0=.a�7��h�Q�0�����q%��� a��q	s�Q�D���	��%L��(5��A6X���LQ6X���j�o]G�&f8��
��Q���� yR����'��ѾI��lL0=�`zEI4[o@�`z\��8���L	���
揣(���IL��0=��d���0������(J6���XN�2�	��5L�o(�Q����(J6�L�k�_S��Xg�����(J6�L��0=��ds��0��x��(J6�L��0=��d�b�0��x��(J6���`zEɦ`�a����Ǉ(�F�α�~����wdv��9@=X|mg�S�a%/X�V1m��S��V�UL�)�T�|����`5q���Sb8�+y�j� /|m�4�p�V���(^��Nu�������3©�,X�+��̆����Á.V0U _��T�|����`�{��>�����{���� ���ԇn0�P��'��A�&�䭟���D_^В�vϼ������%?h��?��F6}�'�AaB7���[?�XZ4Y$o�c�#�!?h�Z{��o�Dd^В��l����ʼ�%?h�?~�2/h�Z{V�o���yAK~��3W~x�iE�Ӓ���L��ˤ���Z�֞���[?q����=�燷~VǼ�%?h�D?���yAK~�ڳ�~x�'.����gD��� �j���>�&t#�\�����E�E�K��)?q����={쇷~�2/h�Z{��o��B�zAK}h!L�F:}�<�V��]�O\���e�O\�-�Ak���᭟��Z�����[?q����͕���~�2/h�Z���o���yAK~���~x�'.����98��V��˼�%?h��uH���˼���i�tD��o������G:������,��>�H�����[O'�<%��i?q���yAK}h!��O\���e^В�6�����˼�%?hm'?���yAK~��\T~x�'.����9���6��yAK~���`~x�'.����9����O\�-�A+.UD��O\�m�fI�۾%�[?qYZD���͝燷��|xJ��g�,���~�2/h�Z���o�d������B��'.��e^В�6�����˼�%?hm�L/����e^В�6ק���˼�%?hm�R/{�"?qYZ4�A��wD�2&��QP�t^� 	�*��Hs�GT���=�#��Ie ��H*y�GR��"6��@��T�[�����^'<�J�A�{w�H*i��8V���^|4��Fz���%�����c�`�w�jձd0<t��X29�ǒH�>��@��Z�����K����T�u�p�4R\�fHq���.ȼ,U�8d)�+Y��C���T�y�"�Q�9^^3��F�urt��R�2�8Jt����d@�F]�7�F�/�c�6Cw�ݓ�k3j��HM:	�2�AfT&Y��Jm|��L#�4��VB$j�8�8Q�S�y�����(�Q�e\y�� ��2�YX�R��k�:�]�*�$(�tA��hX�*��8�����ɑ�D���Vy��|&�ցN�,HK��C��i"�xۢa��D�N''*�mr��N�&'*��er��2LNT�SvɉJ|�,9Q9�0:Q��x�ԝTSeX�uQ�FC�<�U�5�ց�٢��e�G��A�D� X�)�8QQ�n_7��>�2���4�J�%%Y���V�ad��U
�D����A�P9�x]��T������0���K�E��%ZUY�R�0<�"'*'[�D�d��P��Q�j����DFiP	��R�a&�[�D�d����l�.2UGƩs��6?e�(��H�LE�:h'*'[�De�E2��bz��V�ţ��Ɏ�˶r^ݭ���>��`���5"!�p�DH4:�DH4��DH4��DH4���h�B"!Ѹ�D B�qW!�@����ŨH��Ʃm��&��FQ�u&��&��FQ�&��&�GQ� &�'�GQ�U*&��0=��$��gL8�������q%�^&�`��q	��(Jb��������Q��zi�	��%L��(���/&��q��(Jb�����I�M������q%�^u�`��q��(Jb�� �	��L��(ٴ]0L0=�azEɦ��a��q��(J6-nN7)����Q�l�&��0=��dӕ�0�����q%�����!L��(�t0L0=��8��=�Ä[��-o��x��(J��6L��0=��d��0��x��(J�*L�G0=>Di���Αe4���O U򂕼`��qe4U _}`%/XŴsTM�WX�V1�BS��V���]^���������5
�X�V�x�k'c�>���b�I��
�����vRE����+y�*��4Qh�@���J^��=�~?������쇷��.Oa�����^�'�����{����O��-�Ak���᭟�Z������[?Q����=����~"1/h�Z{�o�Dc^В��L����ȼ�%?h��?���yAK~��3>~��e^В�������˼�%?h�+?���"�iI�O\&��e�O\�-�Ak���᭟��Z�֞���[?q����=�臷~�2/h�Z{��o��e^В�������˼�%?h�YW?���yAK~��3�~6&��˼�%?h��c?���yAK~��3�~x�'.����g�����nEO���e�O\���e^В��l����˼�%?hm�?���yAK~��\	~x�'.����9���O\�-�AksW�᭟��Z������[�'.�����D���O\�-�Aks��᭟��Z���v��[?q�����Qㇷ�N�y:J�'.�~�2�'.����9����O\�-�Aks�᭟��Z���p��[?q�����E凷~�2/h�Z�S�oC?q�����懷~�2/h�Z���o��e^В�6W����˼�%?hm�9?���yAK~���y~x�)ˇ�4~��O\��˼�%?hm.C?���yAK~�ڜ�~x�'.�����%���O\�-�Aksdz�m�'.�����>���O\�-�Aks��᭟��ZrC{Ut,c�Yu��@�
�����4yDU��<��@nڑT�Ɏ�2��{$����#���Ie ��H*��GR� =��@��R^��]�:�F~��VK#�C��%���kBǒ�H��e�cɀt0F��n�K#�CwA�%���ǒ�H�н�c�.F��nK�J`�x�Z��d0R<tQ�X2'C^�u�'eP�Ih�I����0�2Ɋ�T���D�d?9Q9)�NTNJ��c]%UD��-�2�y���ª��4'*'��(�T�'A�u�Ӱ�0D�BWY^Ƒ(Ocq���rR^T^�24�	�u��8�Rā��Pdi��4vh���-r��i���D夢r�rRO9Q9�_���TvNTN�Z'*'-��ԝ�2�⺨C��T�J��J��%u.�<�N'*'����C����!�D��p�rz���$��42��4V��q�JA�(r�T;�)*�Ք��}Tɺ�)��tX�AZY�uQ�u(���-r�r�ENTN��u�Q��/�(Hd��Py.Uar�ENTN�ȉ���"Sud��0�i�k�SV�2�TQ�T䩃fp�r�ENT�[������a��z����_.����ٲ���\O�����Ų���~���4q��W���,X.�@͎�/k����AB0$v�} ��ú��+��U�`�.X�Kf�qp~�0�"c�>	.���%��%̡�Μ#�p$��f�QX8!Nx������
!H��C���\�$�)�+b�tN�i�>����-�V��Y�e�!>�c�2~��3�6�P����B�~F�Ϩ>bKe��X�����mxI�4\3;=eծ��p8�s[U��N�xE2��_�b���<�ܕn���	E:ͦ8����C�ʣ-xP��Z��
n�)�v��eY:+�|u\�`���;�8P�-�����b�-�,f0]7b�n��]��gZr��Μ��mɹ󞂋@��h7/;N�@�	�${^����LCҾ���iL�FA���-�r����hS�Yۦ�\7+��u��ҫz���Z�'6���.{lsM5ߕ
����̎���	����a �`2��-�8+e�``}��tl�d�N�����8�	�'8��[���0�q�|`M��kZ�S����z�jvxLQ#�F>V�l�B�Sk��	�|,l�6���x�i�Gg.��0ʠ"p\�aZ�Z~�y��3��j��~Y�]���i6/�v��hP�¿�������~��&| �S'G|��'|@�3(^e�ce� �h� ltߧ9?�A8��'�!*�B����L��� M�3�ˍ�q�� !~N� ՝�A���t�Wp���O�0�:p(ȃ8J�y)N�HC�s�xՁ��
��c�m���Py8"x4L�('���� ��-����G^��8CgTF�``�1J�\r�+0Ł]=�#��:�8��8��8뉙�c�Ā`���w���!�ρE�I����O�b\C��P�Q���gp���(�'L���M!qޔ���S��a��C�=��~q��F�zH�Z��H'���弃À�3.�i L�L1�#A ��:
B�|�=]��|0|��
8Q<�y����"b��j�46zo��q4z[�GS���O�p~��
�~�i�,$�!��H��G�1�ЙR0��	S<D߀�)T��)T�,*�_�*x�*t��b��R�ǆ����^��iw0��1�Q*�`BP�&j�:[�gy�?���af1	�0@ y� @�� ��Y�0H����a7�ߎ�!@�zl8uܴ{z�c$������@b. '�;=�@��g�s�a��0��q�.���i�t��a��� lZ�r۶�a7��܍�6p����z�`7���5���
?#�z/o�=��MF���K��rFrD�΀����fn�&Ñ�y��$��@����Ll	�s>�}P6��Y7�|�9�|���~
"1������W��=w��bz��V�ţ�^W3]-�w����o�
Cz��c6	�R���MB�����M�+>
6	3��(�$���`���х8��X���LPqSW�|PIk+5��R��I4�K�7�5-Z��¢.,��Z��]X�Z�&ɅP�|�,I�=�x��$�����mg��o�*p�ڈ@k�\Xl�K [����P�|���|�65>�[����W�/���k| m+�1���+s| }*��O���67�in$@�ʴ��H��U]����@k�\X �˧�l���3lP�I
Յ�?@5��_,��hj��|�<< @S+����08 �/����|�4�T<_>��|�4��˧ap <_>�f�������PC�+�F�㒏�g����]�-�F�/���m5@��3-�k� �˧�l��� (��|�4�M�| ��/�F�����mC����h6��q �kP�|�^%>�3�)���Ч|Ͷ+>��e��x�y����C��ǹ�����er��������O����G`|b���S`�a��	N���`�a���>������#0>�%������G`|� ����3����K]���'ǝEn,��8zv�`�L����#0>���^c�B#$4��lyvb���`�|`���ˁNT�� 7�!:��İ�:�#$4��e!P���0�Ä�v"�����50`���@'�hq�����1O0� ��谇����݆��!:�#$4B{� �Ct�FHh���z
��a�`��0`��F���%��!|1�Ht#�Q!���>h��0BB#�G��<D�ˀ�=f��!:N#$4B{D�Ct�FHh��;��{���qB��\t���w)It�$�ه��bڷA�w���0�P���0���O0<��-]���Ѐ�0������]��=g�Mg�G�c��q�	��{6� �������n�1!����h�c0BB#���<D�ŀ�=Ԏ�!:�#$4B{ �C��b�	��&@�ŀR���~0�j4zi�����@0`��$%�a鉰�w�2��N�o(AK�i�A�F5ԀR�3�/��G�c0BB#�)M�<D�8`��Fhӱ�y��q�	�Ц�A����{�a��q�	����A����7��!:�#$4B�+	�CtFH=[�&s5*DG1!:��"lq�uH�Ѐm+4K�Y�i�+5!:�	�Q!��؈��l�uw%�S`.�AM�j�	��&pC�Ԁ�M>�a�j�	��&�C�Ԁa�JӎoƼ�8B�8]�@�=G^���9�j�����c�e~�M�}(A#�u�������u�}��ov}U��LF��}܁���1�ߧ~�Fñ�z��c�����xc	p�{��X���c	t2�%�I�;V�qun����Z��u��69�-{�P��dٽ����%��\������{n�"���Z�4�J�܉�8��#�{e�X\]ܽ�i,�.V=BHzGt{^�u�'eP�Ih�I����0�2Ɋ�Tj�s3؀Rq"��Qb�yN�z�� ��5���y�����(�Q�e\y�� ��2�YX�R��h��t]���Re�E\ׁN�"ȳ�P]eyG�<e8}d�;}d���eh>Z�@'q���Qա��4i���!s�D���!k�D�;n������uN�zL���s"�c�,���>`����ԁQ�D��}ϥ>:�Mn{����)�*��:4�O偮�����*MQR�ʣ�Zp��;��@�9��#9�yN�z|��w"�3S1 �N�xJ�%%Y���J��1]��U��+��<�GU����T���GTz%�*�<dl��a�ie��EU֡"��w��~���/B]Fy�i�&
�A%T�KU�E������N����LՑq�\����OY-� $RE!S��GǾ��G�;}��������Y9]-����ţ�.\|ދG?^XG�*A�X����L;֭ݴ��Z�f�q����]hlMc������v7�@�c4
��ڍ2j\3�e�LV6��4���R����do2�7�X�6^����6nۨu#͇.��=W^��N�g�l�9X���7T]��0U�A1u��:���G.r��("�Q��<��G��;QIP*#]����|�4$Ѫ.��<7�T�In��,EՙhZoi�*��6���}EZ��C�z����E�Fj]R�*�U^����yOY���b�S)IZֶ��w��9�VvtN�ߋ�ۼ�cN��C0���F�q}Ykj�u�.8��<��Z5CΝu?,k��}|��P	��OσG����c�C'Ot��=ǈ�Ѱ�Ns�1ϯ�7�v�Eܡ10��^u%,@6�5O��[w�\��l8�l��������W)t�4��_�������{P;AOa�E���v�.B�r�9�x�)��چ������;R!`rj$s�	s�W|�4d~��Y�]4!k98�A3�89Γ���h"�Ҷ�{��4��q��I8h�\�atѤ�h��F��cC3�˂�-4]}(��G��o��*������k#Q�G;��g�ew�qe��e��p(�cǱ�=�Zr���Û���n��;�^��i��G��Ůn������U��jz��յ�nQ���]��XYn���+꾒�W��Jm^��+�~E���2٭M�j��n[�����l���h�.�K���t�.�S�6�nԶ��e[�]�6m^��W�t ���W����Kmq�.ھ��w[��EI���G�-�n���ͻ��n�<궏��C���[Y�]aW�w�g li�t��骧��M�i��6�A����-I٥)�PdO/�2م���z���f�z1��ݮ�uM]����������V��]_�U�jVS?J-;�x�u��y�5�^,7�r5�쪵i�ѩ��l17T^E�L(�0�R��H-"�6BC���g��]�E�N�(Ȓ�8��qz�,� .��IR��淫l^��qZ&��X,gy�v�4ɴh�,��Mk~�i|^j��ҽ?�zu��N�U���Ţ��X<P.�n�D����_��-���[����r�&ݨ	'j*u��b7l�&�3�ۆ�r�F���iE�n3��EN�t�TL9�#Gt^��]�iDo�v�K�[�_�����L\h�؉V�DK��k��dC��؆�u���NMm�ꭴ1Jeez��zq]V���~��go��.�tq�s�*��tq��Ŭl���cm�O@E�:Y���\�qZ�a.�HVM�ꗛ�ŲZ�����������2�� !:a�GePB%�y�FR6�����#�R�af��� �ʅI���1�E\�{6��[�},S�v�
ŕ�����c�\]˲�v�uo�Ϳ�,�oO̷uv}[��7��r�rN��ظ����$	�*�LW���E�:`�W�r�X=���{Tʸ��Jʠ���P)� +�i��a�s�����>���X)UqYW��:�"��8L�X�u�l�����l^V����[�3�����'�����bSz��w[�x�򅒓��w���~����qY.�����t��.��u�#]W�}	����ҁ�YA	�̸cI�QR�C�f�`�
Wj"��A��.��H��*��O��Jd7/�J�d�q�R�	�T*�sU�ɠ�e&D�CR�v�T*��bPeIiV'E]��V����_f�����&�������J����駟��/���~��~��e5�],o�o��zY-�u��-.�z�z�¾+�z6�&���7����	��^Y�����{��߾��|��o����x������^>�~�'_|1��U��ue~�������6{{s]�N��;�m�O�>��ޣh5������~��|��;K�z;[��g�ۉ��Z.���r��:)g�g��zrc��C2k,d����r�Ҿ��Ę}ϵ	����&n�{�8��yl���牉������铿=���~���|51�M���?��.���ܮ&�颮o��c��^<پ0�}��lnB��z�ߦ&���T��ּ��Y#�/V���_7�����������{����>}��뗯,�{A���ji�4Ҳ'R��v���g�{�LW�5��w엓Ė��(2��"��̌���
��2c�ƨ�7Ƣu�6���Ɗ�	1��y�Z�3�����fo�I6�W�'����H��p�*��4�v3Y-�Ho�X
�I^ݗ�dHe��jh��-f�d1�j[h��{L~}�p�):�����6�˧ooV���^X^4z�M���������?�1�t�y��?lIN&�z�`�g�&_~9��]_߬���&��F�n��~�য়~����7�<y��_M��ÖK#We�˗�Z����F�Mf��#hxflC�^�z9�uq�0��R� 83#w��]\<���\=ڧb������Ͼ����=����I}������r�+�e�=�=�_f2�߿~���˂m��Z�&�z���R��B�Ҡ��|σ��?����X����U1�]-<��Cx������tV��+k~,�
�~���6�޿눖u�_ۉ����~h�]�mE�~|/9�L��?؃�/C{��AX�]�����T`���ark���ofa|X��̀�zv[�S[ {#
;��+1�ʽ�L����a����Pn��}c����͛�����V�����ͨ�oC'��`������Ͽ������?����'��0o��Q������������A������j�bk�>��>�����7�Xg��f�G���΋wֈ������׻��Vt+�/sc�[bk�Ք������w?�W{�l�vvqk'_\N��|f5N�n���}j��e�ǚ��.��ůoo.'�ۛ����MUY�J��i3�1���lU��õИ�[��w�jm׎B��8W���כ�q�"n����ڌ�����?��W���.��������z��p��h��x�����/�p�&���~}`���ΐ��b�ݎƭ�����J�>�bn����Yf���1a���jow�ڈ{n�����~x�6%cWwK+�Mx�o��k���������h��Xۡ1�[7f�<�c9[����g���������W�p��~664�f8�+������>���W�/6/�<�7N�@ 0y`������Tr !�ԿOH4�����@�ޛ��+�������l���Z��=��{k�t�"��MM������P��֞�0��a�.��Uy�ߎq����x����5C�d��wq�����l�f�[�5��l�߁ �����I3�o'o����r��M5߆\��S�b��F؛���z�'�;�%���_�|kU��F����jS��|nۃ����[��~<�x�6��7�v�j��h[�g{�_��{��CO�J��F�m���MP�ϑ�M��o�h�N�09ʂ/䶥,د�ao	�GkW�l컙���l�١��p��S�|3���w�~x��>Ѽz=�? �G{�`c/���M n�ƛ��yrS��=���Ϟg���i���޶LԮ7��b�̦%;Wo�V�=�]-�b5�L�쫮��x ���o�d��ۅi]ݮle�(n]�Z�Ɲ���]KwFt��2�I.�&�̶��(�F�]�y���%��֢���&�$gF�=�|p9�3m��~c~��}n��]=5�6T:~�h+�ۏ�\g���g+6�m�*�6ٚ��lb!\W_�(^���4���?�>h�x�����5A�a�iy��wܫ��v���x�﬩ܼ��?\�?YZ�?_|�_v�Ǌَ���1����]^����Hɴ\��UJĥ�������[�'�����6��ƌ6Q-*c{o�]�q����=�~�yK�/w��*a��ԶQ6(ٹ���3���ы�ޖ�����[j�X�Z��7_ܘ
I\�c����Ů��R��R�L�g�:�K���6����d�!&�M��l����5�a/�YOi�5a���&1O��G�#ݧ�7�w��<���>]n>�I��R��i"�p?�_#2����?&A�'��7˾Z��jY�ֲ�e�ظn�ԍj��gv��n'���Qj��k-�չF�f�������hS��H�y:7A���� yg4�w'����6��;����ٮ��/����=��cu��c��X��rr�d�"������ɮ�6�?,�S���D�Fs^6�m�Fol�?h�YU����,���&�X��1��O#>�m봈���M�o>��w+t,�a�����nf�6K�.���z1������*��H�4
cG"I/C2�Vq��ȼ�^5[�~��^������&�Y�s�+��.O��
"��"���,�_�$����Yp���j�:*���R�N������d�R���V-���Zw7��ZA�w�Z���{�?��N��.u��%x[/����?�Q�����a��ޮ�����ˋF��ߤN�>�;�,���O���|��!�]\�0.����Y~]�-������v+<o��]��?���j�/v�կƕ�W (-�J��J�a�嚽��*}�(�����``UR�e�:�#�q�"�I\�u�J��T9e�q��D�w�5������W��8L�[S����ϟDf����&[���9\0tx�)wN��f�����i��N.t�LGU��Zib�Xe��e�8YR��-N��r�X��h���&!��P�ۑR�k�P�D:�-F-%%=��:�^��)\c'u�ѕ��Ȩ�}�
eJ�´��R�)*�@���Pg$j��%ER��������6TWFA$�ּ��el����J�ٴ����^������Uz�{��>:�>�:�=��^�޻�z��;3>�$��VX����\��8CR�D�A�y���P�AE��0�<��c�)!���j�!_J
�[�/������Ѱͣ��Q�)o4���x]���t]���:�ޅ�Ds��S���2��w���ټ���T�xgIZ.�Ư��f����HT�u��b���ʨ4.���:I� uaD(4z�����hm�r.Β�;�M(�;�mݎ$4j{� w�x���{����&3n���v���{Ks=+���n��n\�)�/��/~�D@M��Ny�AN�%]t��k����F�lO���О�	��͊�%%�\IqJ(�d��ak��V���Z+���.ݖ��ͯ׋�fM��;R�=ܾG~�hW�ޓM6��Q�8��򢾞�|�=�bV�c�z�bWw�Ac�'�^�]rM�@݃i��o���͟�����MV����m�]5t��=�?������=��^�W/g�]�Rݽ��(NR�t Fwf�,'�U��k?�J�8�C���@�KJ�+2�(E���:��	�:�v^�(���\��&QADu�iGR�����H�hñ���} �>?�@�U'��Z�ad�zy%�$JCE��i�PtJ����ݐ�#;�������{L�(4CQRL�ҌH�^EJ�85^��8a�F�l��р|rW�<�j1g�T�;��ɏ;$#�04�qDa*�Ȯ嫫DƤR�5a�H�[#�#�f��2Ќ���ƾ����6��$6�.��`�������\�i
Ɖ�kcmK����7�J���B�lF�_:��zP�ak�o���.�Ћe�Z���Y�����6��o�������o�(n��v-�H�o��})�����<J�펌��2{�	��{�Cw������4�~�[�m2�����e�{����~���)�V����
��usx����J���/{��[���b/��^1}�ث?]|0�y(ji%DR!EM�DM�EM@EM!D-��3>��Ab�A���J��O��p�]AsD8�7Ҹ����A;Vx�A�����b�D;��?��y��c։{X*NX+Z�TY}�B��T�_�%<�bg��s�f
P窦St�7����������S?��u�5l�e�&*s,�B73��8^���:������#��p���~s�a�+��i�]ҹT�.������B�+���Q�U\G�D�Ӱ�*ϴ�#�"���Xa=��9$��R���{X*>C�R��0�g�RI��˳JuDz-��9�"7�?jx�����܇�����w��8̸;���z��C���0��c)��Vf�u-�(���
���b���)F`E�a\��[Cի�;��smaut�:֙B7�\���mz�e�S��YXG��.AIK��:��?(��Rg��s�=�N���A�%;ME�ٶ>�c'V�5��O���}©{1,V>�THS^�S!�S�E�U8�z�ͽX;2D@z~$��\v��3��u7��� �����v�>-�TZWQ�+o}�G�@���G(�h����=�>�cU��?��/��ǝK��u����}�Ǯ�9���3�e����#�}S��{��ݢ@_�)� ����4�=�~�����z�U쓎����G�1��{���~�������~!tB�9�{�}z�����0?<��	��eC����!�+����[�����A�Ra���7�.���~r��<6�8����X1K���i�A�Ԁ ű����:k�kJ�(�.feEH1;f���2/�bC�lo��i'1�Nb����T�����R�b��:O%R̎m�.b��i�6�����h�NF3u2��%���M��^�R�bW�,�bvlFvl?F`1s^�o�nm�.�/@�ey�RQڿ��(�*fyY����c3�c�1�ى�p��+f�E��K�t�f�R�l��Z���q\J��YFu�z��m�:P�4X̜ϔ��7V̔�6SN�L9i��R1�[<�.����y��R�"+D]�	Rdݎ���Ĉ��#��D���s�)�E6tҌ��flm��G�b�v�at��,-+Dl�,z30<�����74X�������n�h��/��B�J�~�
[g�JE���幺�v���>��6$�0K�[�C���c7|H�5M����#PN��������h�<j��)ƀ�=7�yX,��Q���[��i�)��,�=�h���p�q��ga.������������NTiB%��9�&ưIhEs���$r16Nv�U��Xa;~v*�<��U~|f��W�O�[�/q'O��u�N�d����O����N��sJ�OB��Kjn��vl�T�u8�:�$�0��g	�hp���5��	�v�S�u��CF�3Nƺ�?�Ӧ'g�'c#��س��[��Г���\��(�[�ci��i�s�Q���"���O��r��r� �"6rWJ�u,5��f��]_?���Vͽ޷����6����*���w�����g���m���PK   �WWMYMVx�  d�  /   images/010d914f-59de-439a-af91-012b754a10f1.png @翉PNG

   IHDR  |   >   ( �   sRGB ���   gAMA  ���a   	pHYs  t  t�fx  ��IDATx^���]Wy�?��ۛ�U�e[�r��6���C�B�?�ɤL&���!mR&�@ �0:�ƽ7ɲd���^�^N���YW6a���������}�^{��<��#^��R���o>�	�^~E�������k�O�Nԥ��\.7y�n��5�^U���w�w=?.ߦ�ȹ�~�����忾W��>���k����{�9'������u�������e�������z�p�~PV��嶿�jS��V��^>?J�?�z�:���������ݽ~�]~��:��l�����~���a����������.�������k�����}�H�_���}�_���~�������N�����[��a��7��D~�y߳�W ��i*
�u�-5�u�e��N t�f��!�i����A�_��C/�>p�x�GB#����z�w��kp���/���V�>?�\�����K�p�/�����xh;�ÿse���;�#-����p��/����+u���aa�������z��x�6ľ�\��_�s���;��e�\/���'^9��gР�Z>��7w�>�_���z��e���_�&vj[|�<�~߫�~~��_�5�����=���]��^?���}}��_�;������"?@~�wm�a��Â������r;�������A����z��s|����m����6��~���~����
�7�h��~������T*��A�7#��OmGh�����Z1Ub��Usm��IΩP��GiÔc%@���	ͧ��p~̕��F6�tw���K�^�x"��vb���3��ϗ�h�A�M���l�OQ�۠㚶}=u�p�oE��w�uʠ�V��+�;�����G�S�\�� q:�DF�D;U~O*�ɪ��*��k0�kj�.�S�E�C�^.�(��~+�өL\ժ�5@-�N�k(,B��uvP�N�\�}��D���zI+����+J�!"��mDT�%����VC�es<a�l6�[��o�*����6btŹЧ����m�v� Ӧ�hK�UoF�dUk�KmpM�m��A��0�R9�SaF�M�}?�<�jCv}\�B־���h4���Ru�٧
UI�	��	<d��:�=��;�$���D.�vB�p[mOܔ/���(8��I������S_�|g�M�K�M�V��]J$�ȗs�a���9�l���Վ���V����I�z�c�S�v����>��$���.mt��\�u�e�VX׮�k�u-�g� ��r=e��H��G�`q>�\�6�}ۦfR\_�h��c�$�-�ѧ�#iᚴ�R2ԡF�]6o�r����r�)�ǌ��Q�*�HQ︚��2��/�ﴨѬ�ȃ7���=�P�:ڷ:!��*�$T�����~)+n��Qd�*�r~
9Wp�2mr8	�4j��G���r�_р4 �\�8���l�C����V�}��jSY���f��'���TO��J!�f4I}���~U���eZ�����Ue�i�Ɗ��r��Yj��o�Ҫ%�+nV�����c���+�o6_==����'�|��N� -���� �ƭ����6��V���E�P}��֤� �<�vu�Iœ�:�	@!��XS�Q��*����"���K�84Ɔ�k;�3
��ATv�8�~�F��ܬM]���ϴQ\$(\��
����F;TU�؜�/3��e��{5U��D�g��p�� � �� |<��]������r��8 ��Dى��u�E�#���+�'Ǜ�2��/��ڇ�!82����à��͘,����F��-��5m"�f0��F>)#�P�猋��NUL2��"Kdj�oQf���z�o�2\ S��c!hِ-A�GB��N��&��,`��.��C��+�#�� M�/��*&	u� �-�$�� � ����b�'�Q�P���|���v
�L����8�uT����p�<'O/� �x�ղ}���]w�>g�>ϒh�!���/���q{����}���SoO�gg!
q�_W���IeAY>^� ��mᕬ�w O.�_f̼�ϙ���A�%�:�%�y>+��_����.s��� K�?K�st��$�H%T������Jc���"v�rQ"��G�QT;Ax����s��M_B_�-�B}���q+��|�}0A��Z�����c��-L!�4b_p�8�kc Z�zG!-�8ފ��g��Eku�XTi7�\�P�=��Z��k�B��o�ǒ|6�ޖ����lq�l�..���(�ͫT�r�AҌL��p�6uI�H���aE|;�]F i��!���mG�I�Ag�h �{����X�Ar�&B�3��TU]����ߧ�_�ui*g-�^�����������'U�qv���J6�!lQy�`������!� ~���xq\G$���uΘۀKz�C�Y �W�F|0��F��V���W�/7(j��)�c�a����gZqn�˩���R�����H쨼8���eP"P=N��n���9��a���4�Y����jY�ͤ)�X�K�ap-���M��u��p�2kM���РLwT�ٸN����w�rOBA������7
m�a�@|�yU�dV��y��u�ؙ�w9ӈQ�Y�����G�q��U�vT���4����3���E6!T�ZJr�g�|�"��7�=ѐ��t�o� ����b��Z~7Hف}��N��E�����7�*v#XԹšc�A�Y�m���q�_Keԃ� ����0Ͷ�D�nZ8��ef�ܽGx�3�P�e�Y~����W�����9�n������8[L7��fN/r���&�}�s��8��t��P�(����WӸ(��Ӗ�kb�6m�x�~w}B���-���A�*�ڹ���^n�[D��n�	-�-g�}���:��RUiʠH��8�A��l���\ب�=)���R�A���F��3�u4@�{�X~9�q{�V��9�l���F�Ͼ�2�uel	ٱ��I�n,r�m�U���u�`��D�:�q�&g��d�7E����G�g�1�*�V�s�ud��)ײ�rF���@�RW�j��yև�IR沬�/���Y?�uY&i.]��٘P$�(�H�؈m����Q�U�!�%S���v3�Խ
q2���-��lk�Y�;�d�wi�7�:�gW�^����]<rHſ�#u>�ղ��U%8�ҝf�0�m�7�D��J��%"�O�ԛ��}����@|�_G���V^�JK��L�J�� b@o,1����c�v�c���w�pk�)u�,�"hc�l_K%�l�f�ˌG�t�heB]��7�?'��z�iSJ�?���	FA qH]?�؊����)ݙX1����&Q\h��@ lahu�̬98woc�����m6�m����(k��U���h0�R�2l����Xxl�M�W��%��*�z�'��~�f=�wR��ҷ�������8E����P~K��i%�ڷC�Z8I r]l�,W5̆es��:{� 4��v+���x@6k$V�@�u�|��mӤ>K��}����V���+42�J����k�)��~�Z���|N+�����BU�BC�`��I�C��� ���J�m��.Б��9�W�G\OypR8���m�&~�~��9�6��xZ*`3o��V���?�]f�&,^��nR��.� ����9��^�e�,;t��s}(㵌*|���-ض�����)6\�2B�+�YE��$d���F�[_/wt�k���CGt��i�����;�u��(iw�H#������Y/����!��b��B��f@
�	�C�y��2��@=}>��n��������
�a�p���4��e}���^2��q�l2e��l԰�w7S:�R̨��\/j�:�I5�/�v �\�;���R/]�žɲ^�X��a;p0p}M��3����e�\����
�s|��ĝ<�}|���7�P�Vx'�6!=�x:ؿIm�:K|��n�FJ�6^���)�b*bݻ�+E%2��������BW3���W�?��3���Y՟{T�}�Hqpe���뚳�K�QD�� �*)���>-�Zzv�!R���ʪ׈H�]P3��dt���*V�U-&��Y�*��9u$�p�T9V����^2e��]�
(��ЊH�[�e��ǺX�4o�!_[E�Mʮ"�*������a`�zD�RT��t�pI������,W/p�]_(.(���՝ך5c��^ІNU;���Gڇ�BFC���/���b�`�
�b0�p�����	�FB�ъ�8n���@k���8h����t������)�@ ��!|�;�"N<~|F3S��՛��Yd��$��6�_K@ð���^R��	������]_�҆Χ�,t�0����%)�]'!��΢��Ǩ#e9oN #�jۛ��(*g9N) �l���E�//�K/л���^�N=��Z5�
�,tjx�����B���Ö� h��	z��&���d*8�Sek(I}��Ln9kpʿ�� ����ɱ8���$)��;w�8�`�Lɤ��nx:��S�>t�j��n}כ4ufZǎ��f�k��pR�a�*�:ߐO�2-���$������oi��\�{���A�9��p,K���MY�K"�L����\�ci�kI�)�?w<٢m��p�__��*r�����՚�闧�*!�,Ӏ�l5424��J��=d�5�j[�P��e��޽��4�t�\�4mHc/Y��X�v�8��{���F9�y�s�w����2��Mt(���v���1�c0U}9ӥ�	���u�F�����;ioTgN�T�Z{j|V�֦�97��P*��t��'��������m�?]/�鲜�s/���X�]���~y����`�9���ۿ9�̢�^��G��c�y�#��@�c�z"٣�'����_��_����O)ݕ҉Sg4?WQ�R�J��YBz8;:/Z
��H5cv�voD�]p���&1�՛�{�k�g�����7��g��|�A->F�<�PC�	zU]�V3xA��WKTf��k5��w�O>�%X�DaNg&&1�/�I���;��POR�V����ER�U��Tk��Fs��� ��\N�ل�}y��*�* zVRU)���D��m�jo~������� �T<��K����w�8��Z���xe,�Z\�������R*������]o�7NMi|qZ������\�$Q8	x$� ����>�g
��k]o�.�|+��
��T�+wɅJ,UU�\�J'UX,���@��Q���9q�^X�(u�G�]��F1�itrp��siiŘ�{b*�{5��i1�: ���[t�3{5[kjjjNS�du��i ��c��lZ[�oVavV����V��׫�f�{�5��h}-9"�Z�.��Hk	�p�RA����Ř�;_�3���0���ڽy��''U���
6�	�qۙ�hp�Kv4��ŉc�FU���d1��{�9������6�Ē�����m�6M�,�S���.t�Qu��|�H�HК��Dȵ��f�U��T�4x���E�R������Xh4Ui�ɴ:���"�OƲ�F&gA������қUg�F����͚��f�o�Q�:uJӳs�����o�6�ztX��#:�~�5���ƙV�{@b ��(v���:u5�u�����(���J=C�t�:�h�/g	~��<�Jղ�)���4�R��W�q�=�ʀ�4mX�C����H����Z�/��LA�>����{����u�`Kh��5*B.���]d�K})�!�s� L��Y�75���n�ay���#�r��7��*z�C~����e�CG�54���!8��&h��,�j��I6x��շ��"���_�l�?�c�|�E����47�����oܠd�݂۫E2Q=��N�����9YD�%0o����U9����JEs��y��$Zr�e�/������p�Z9���n��z�,&!s%�j�vǹ&�!��<���������;z4d(��9��m�>{!z?]6��j-M��)��S�"&8���躍ʾ�p:�(y��
��`�-<t���`(]Qeda��fY���k�>��'N��m��n�6��GԻ�&}���	0j��TT*0,���ȼ1���p]�]ZT�Xҕw]��C�C���;��
�6���JC�����9���ם��շ���j�-��?���.Rl�*�x� ��ɟ��G���� �x�Όu1A������~X�k�ЎwޡMw�Q��C_���ɥR`�N�--�п"'L�f��Yʝ�+i�E�tӯ��֬��;��6��I95�Q��m,GP��U08��Lk��ڴ�4��D�S K��k"FxM�\3�@g�6������^�C�Eu_v�Fn�T����(�q�>��Qq��� �I����L���#�q;�E���>�m�~����U>�RM�ؠD����q�0��lk ��՗k<�Ж��z|��G��є��z�^L�5�ߣ�ݢc��(v�Uʟ�V�v�\�\R��oU碋�%h�\�Q���ߩg���g��!g>3X.���b�ё�����h����j��Y�]��t�M�Q���ܾN��6��r�Z{������ �]���.���$���&A�C�J۷�y�E�I]�
�
�J0���HBK��M�;T�t���ۡ�~�?hÇ~Z_�������yU�N�\
}�N퓩t�93�t�䓓S��Z��g��jo� ;���촶a���=Y��)�Z�ٸR��������v������=؈��X�S���+�^�h ���(I���=���@�w^�2 ?�q��iL[n�.�˿��ڢ���d��
����+��3q��,�o3�n�_h�duw�ß*A�~����봸z��[v*���B?�Ű�&��'8;�'�X& �8��n"�5��a�]�F�I/�-��u���T:���*=9]���vޘ?:��bY�KK�q}��_�W��UU�5�2y�4E;�h�VM�55��[nTr�VퟞT�YZ9��ͫ�yd6XV�!�Y|��W����ޑ����v�!Z�u���VF���ڟ�K{���R����t�1$���t�+���d�#���a�����^�K��면�yD�<��ΎOBL����z��Z�j��L����*]��RdM�j�NcE�
}+�#[LC�j��3
݅���Ɗ��}�B�V �s/�q�唛�t �7u��]��iu_u��6�Ֆ�ߦ�\A�\s����C�Q#I[����� &E�T���8Xg��;�q�Io���]P�ONh�ڭ��:�ў�K�NXR��굚{��`Js�z�M�F>۲Sۘ0�tΌ�'���y`�V�g�4�ue�Q[�z��46�֊�.M�4���J��"��}����:/�9%r����l�S����� 聍}���J�\R{rIq2�|�ĪYUbn��4�3u�*bT'+%@��d�+�[�k��%�U�Q���4&�1�0ػXS���ڵq)_M�GFu��tp�j�H��
��in�;"uw�� 1��!8�)kV���=H;F5|�fu��I�rJ��ާ��O�'%{�&a4� 鋯V�2A���&���)��WF��F�-[TٲM�'_P��8�,����W�}�We ax�f��{YM�:�����4Y���VMSF����N*��{�Ȏ���7+һA����=�O��~7�&U!P��2�TG��gb�?�����h��+uf�Q]�+?��~\Q�53�np��������C���Q-������\i]�+�~��|�p/�b�vf`p$!$-����ݵC����-��}�Tx�Qu�Iױ�v��� ��w�����ܧ5ҳ���х�6Ø�AժZ�	�۴E'V>�je��iTG�isG9�+�����w�v�F����:w�,���G ]�G� �x��d?a�r�S� ��]��HtіA]���&{ݬ3�ң>�����Z9UR��jlDm �!�Q)+��.����(~���&j�(���P��Q6�$صPd'�B���Gu��n�����V��M>�5u?���+U������x��c
����z�����V/ެ�k�Wm�Z:;���s�hY:�M[!�"��;���ݭn�~�����MT.�}����*�٦2�<��b�N��ښ��igZ�~��T�R𬮾�;U���U��1���\�P��n�n�'0��-�Zs�����T^������2���� Dp�>���S��m�p�����>E/��xL�| ̿��6��;�T*)�cG��[��պ灧��>�s�ܻ?����sT��/)�ç�/�{��{`$�"�|��EU��?��>�~�[�����"�~MN� �u���n"K��V��!�9}���w�ܽ�����k��O���҉�vS�N	˕�##X��=m�xA�'H�{�4sbR�^8�_��ú�'?B�T�Hg���o�%�<��`D�4�����<�/��V}���P�d��<��Ȫ���I�#J�yDӞ���Xc�WHSk�n��%�l��׍��4:8���˃&p>�wL��Ns�c��?�G���K��������?P4GP¸{���wPqFb�����P'g�5["�淧~����y�Ɵ<�:������ c����I屇���P��t�i�����S��:5���?�3�����j�T�K��.D�ꅡ��U���P�k���F��}�}��Rˆ���U=L5]��mp��J��KK������?�SM�3[P6��ƍ��X�$�����8�Q�b�I���A��Zm��գK����O}C�����Z�۴3W_V��]��P�j���U ��}���_�ŧ�'P�l�.��A7����vaŞ��1�'���bbN�_��N�Z��<��M+Z�V��%��
K_��W�i�{߯�����8� �ب�v�J��.��b�%I[W_w������Z�n�D���w�r���r��"�NN{�z����k��_��҉���E�l3β������GPZ}�E5�����O��u"�0շ۶N��l�Y��j&�׳��v���J�WU2�$�R�"�PW_��Gޯ7ߥ����yO���R������em�v�.�y�.��B\Jp;��N���ʥ*�Y���a��x���j�!"z��!d�!ǵ�l)�\��e4��Wk7�V�7��ŢV���X��d�V��z�_p�z��ZSKs�����Bp��5��4����u����;ބ��Ij����~W�/�	�kժu�޾YKSs���L���UW;K��qƃ}���8��Y��a�<%5�]!�k6���߮]��M����$�;�"s�+���;��2����W�t,����O=���=��_ ���Z�)��.�8��?���AT4uv\Í���>H��Dq�?��ȕ��b8�4��l4��=�y���֧�����w���t�~N��\l�T�'h4}��J/����O�DK7wgu=Fr�`��a�3Ͽ���q�]���y͟=�i=��83�Y���~�cz��'����Ua��մ��~փ�dz8�����I��7!�C���h�r�5_?Q�h�9�g�X��	]~�������f0�Ylo
9,]�x�:y��J�g�c��ʡ�3���>~|Q�d5�n�(�3jN�x'�1���f�:S�g��o�L�U�*�;uB��������ֵv�r:���4�S'2�^K�ZJW�Ϊ@���)/r��oC�7oV��N�s8�D2��/i!��s���N��WՅ��n�[���tQ_Z���� m\<xL�jI�������� 7�~�z+Oh��)�L_�����?�j�<�T̃��;@1��=��u�f�������C �-�o�".>rB��~2����Lg��ߪԾc��q�j�Iu2!k۶����:��(0��k��wj��Z�q��¦OO��L��i�����j����?�I�H�?�7�ѡǟ��x]SY��'�,��@Z����w�`.G6`F=*�Oe�r~Vz�>=����y�/����q7*���x�Z@��dy���*L���RK��Q�Q" ,h2P	�kh bS(c�{�gt�,�}᠖jql(�/V[X�e7���������]#����C�&;df�Id����n�b;�5����I?�]=��nu]x��+1��^Vbד_�'/DFZnX/�P���|�m��b�W�5v�F��x�~��4q�����
Nh���kk�|	]������'�شMIl���~��?����u�gu�����\����"{�D
�G�QP��,"���Wu�+_W��_�z�&���'N��ȣj��P��b����\���ٟb%� R�33j-W�TT�XT�P�.ܹM�����O��~-���fE�����^x���^����_�����_R則t����u	������mqO@�w7ty������<��}��܉i]��۱ �С}ʿ��RD9$�6 e5�F���	S��=g��ʴL,�}F����U|�1@��/]��� �*B-d�PR�h[͂WJ�p��S0��ff�8K����p����0G���HUJ�h>���EE�d�߉��hB��a����.�}�1j���ӎ��j���NE�g��Rc &��IgP��:��'�I7�{`���2�KD��
����>@���T�a�$�F��,*�8�!�Uk�Y��rAW���O�	�8ɽ;i�7�Ue��9�~��z�yۻ4�¸fO�+ۣ\W����OT����kZ?�t%�|���ÀC˭���3��c� wZ�0��F�mUy�M h��k��qİTt_^Y t������0���;7����ղ��)�Wԕ';��6u��S��K�$9�	�����IR��T���I�	01 ���^��½PJ0k���#�ֽ8=O��:��*�UB�_\�ť�`�El⦛^��~�~%�0o��16Q g����O��a�	5z� 0|�y�\I����;��d�-��%j= {�d�7��,�e��Q)Uj���r�:�<��G�Q�m��"5-ub�l�챗T/��t�� �����xW���ޱAi���=�������9���m��UIw��%]�j��b�0�$,}�����k���:d�N�Cf��1=<���);*�#8z�����2���òWl?O@��|����S����Q�������`L��j����Q�qz[Zҝ�ܦg_اc���*i��?N�� q^���{����U��U��7�B;.�B���AG��ܽ_e����B�8|ـ�9=��E���{�c�6kh@śo�~��Y�F�OF�g_�x��,:��W���)�OM�VZP��[=������;�J�����Y�ɹ|��.FyU��.e�0����.��*h` ��L�zW�Q���o��_����=�f7n`+ m�k��ٽtjiF֯W/���=�X��Vi������s`�` U1���TyQU2: � �C��S�P�V�x-�K���D�'��� �؈;����ְ�������׮��8�o��_���2����%>��0�ġ�k���R�/��/}=`������ �K���������<�e���g5�({�Q5 �gO#�l�4h@�C�����X%�§H��5�<?�}kpP {�ŗj��i-��z7i�v�|���a6�$���D:I6 ��o�F������|n�?t9�G!E�o�G���T�vB�j�`E���M@����il��QԔ��<�S�\��]Qvo/�����Μ���Z%�J' v��Z����y���&/ؠ�nPe���[ǈ;iUkE����7���?i1^��y=��%�a�Vh� S&xG�&� ��RME-yˆ�p�j�I�3�~5�J!+�4L���ګ���qq�O}�N/lg�����H���2p�n@R%Hf�C�E�����u��zu��`�	s��n�en��L8��׼|=��V��[�U�,��B��j�%�k��"���%V����yd`�˪���o.┝6{o�)�rk�EL*��&���5a�w{�87��w~p�Ab�1�繾
MNy�!�����&l�-�˧�Ë�2a"�C]=z����k��W4<8�?�����?Ѓ��Szرa��L��ͭ:ot��*JPL s/�
���x>�l�L�E8x#g�^�b���윍��=��V=˦A9豄n�do@#�_��okdt|�,��;�����Q�?��N�lco�2�Cjr�.ŗ����zA#�[P�"���VȪ��٨g�<<ث�����#�V�ک�v�=�
[ HR|�K�r�z^}�z�~J����4dm=�s%�[��D!��bqA����3��k�.�|��z��Gt�Ci���V�\LX��1���V�4�ݘ(Y����0�"��^��I���c,�ے�<�C�m�wK�k����o{vR̤� ���G ��6��l��B4l>̭�S*-Q�ZS߀��wA���ѷ�M�Xw����/_��\a9㍦Ԭ�5
Y�.�o��ݴ��ߧ�[TbHY��k�YX�y崳����Z��oc������-��^���
Ǹ�c�
�>���d�]D$����aY��*���S!�!'a|IX�?s���ad)@��{�/.��<q�P��U�D�|F�3��܆����u�4����o�w�$^\�<w'y��6umx����R�����!�3X:�hdh���b\�7�χw6�S,r��H 5��nQv!�f�Y�4�MZ�x����SmdD1�Α�cZ�YБ�{u���ܳG�-;��l��ߴS���L�v��	�m�N��*��:���!��ۤ�2?fho2�õJU���㺘4��:�L&�s�Y�� �H)W�H:Y�Mà��5�\�0 �.ȵۋl�؛d��Aӟ��]/a8Aa?�G@!!3�'z x��Tc]d	0�X:��4{�Kd]޷�3d��4`�w2̔����	@��X$��尕�rl�n�����J��5��g�8�=y�
PlQ?�y�YX<fW�V�I��ߝrG�S4�T��2��"�B�V��$�Ǔ����~��@�O�VOO2��lCٜ֯Z����k���_�^zِ�����G��n���{��y�,[yH����nJ�!J���p|FF����3��}��W�����/�A��`�5Z�M���է>�Y�93�$eY�������Y�\�2�6	%�a�,�Ys�聠!��;���"�#Q�h��n�N7����{�$���=&g�ZL]���Z�;����"-C��lԤ��#��DJJաSȽFV�.��V�	������������w��� �<���n�X޴b��x�8���p�E2j�.@*�?�{��ѥ�n܃��u$tYc��8���6 +!�U����E�� �{�P���}��^Jd�U��ԏ:���I�Z�̶�O~�t��)]u�u:��-���7����܂Oc��_�L�rI-�4:�g���I)l�U�����.���e���nEpr����-��3�RPa�Y� ˙�*D���a^|9�H ;l��2�N-��!�.�x��B����V)�v����0���R�{�@�(�3
��\\ct7���(�Mر���y1�";e����~���p��<�t/�%H=�Ѳk��������l��A����W'uW����o�JJm�$�68$�0i��EU�]�\�/�p�%EǆB��02���cꯡ���j�~ȿn<7>qZ�Ds�R��V���)�ے��Ic=ݫ����SƑ�K�*�yi��k(�w�k�?���hV�1`�d��*W �ixʚũO�Fٌ����Fd(�O3�`�����Q̬`�Q�Ey�3�m��ة��Y��)��Ld���:i��е�8��*I�l'Y�\w����
�f�:�7(���<��*����ؠ�q�X	�G&����Y�^��)��*�H�ڈ?JH��yʊ��uvת� ��Ҭ0�O���0&�W��B
9svV�%ڇ\� h��-L���:�
>���wQt����qmo�[iH��ڶ��ma��Λ���#�蒀�?q8�'�tV���oY�f!, JQ�E2�:��l�ؚ	�C����{��eH���,?���Ly%��IBeȀ�2�Ϲ&�,ؘǐJ(��*�L��̪{�Cg��/Z#�ײa��h���i����@�Hs]�ֱ��e�����&irr���w��m�����s�WOowXտz�*�^�p�P�ܫ�4ъW[P'2���8^1q!��tl n�Vu�6"*|��� �:�������������S##0O��QfO;�2�U�8�L��������z�GC�Y6ץ$shh0`�mϛ���Y{y���cy\
'@dћ1�۩��~�y���ʠ�_�S'U}�>�l�п�I��\�E������6(r����J�����e���>�u�_�C�N�V�s�e���զ�6���?�߭����*+����ר�e���a��E��b����Hd���`%9��ǁ�l{�S�"���;�}J����� �׭���]ݗ]!]�E뮼X��ƿ�����>��Z5��+A��P�������>)7��5��?�x��������|�7lQc�&uN�����+��@�c5r�.Re�H����w�P��- p��ch�1����4��4��a�`;��a�/}X����I ImZ�����i�r��>�sy�+�e���f�Xa�#��
��8[C��/k�W��Ud�vE({z������b�6;SB���sٽ�w��5�,xar�^ap�?�zޜù6B�02�4pV6�U�+TڸQ������hp�5��7W�`s����O�a�����=���������V��j=�w��^��a.�!=5I}�-�3.���%�u���������s�g)~O*���~��{��J��tiQ"E�T<-�^�G5��wi&��� �Lp|��'m��_�C��թ�y���Ĥu':��R_��m(������6�X��~�Gt���1��+�ڶE�]J�8m"��9�@g� Hв�N� �&9^�������\�LW�<9�8��#�Ħu���uVY9�Fw�V]x�^����zw�����E�� 8�+��\Bf��: ��"7&p���?��h�N�ٯ������`F}�4A�1��.��\'���Уa@��Z��npn���dxi���d���P_���p�>6�Z~@�l^S���U��վJ%L��X�ø7L��;�S�`"3�b���#)�jv�p��,߭�8��ϲsn���dљ�7h�.<�����MƜ�0��p/�?0�|��-�tAN�6��R����j�[_�����<�;#�����&�K4��@*�4��Mw�C����>�
���1����L*MEj�Ё�X�?���
����&Թ�^���bt��s�
�P��������:���]�I��z�����o~�K�$8tW���	xQ���'cޟ����z�-7h��j��Zw���v>���?���e��k-u�430�񞴦ʀ	B]�B҃����������k2�QW�W�E�`X~�����7h��k���M�ӱ�Ӻ�kw���)��!"������s6�~Ҵ=�8��`�m�ڡ��oS,}L7��V��w	DlDKKsJ�yA�����C!���_P�4r�������_�N��`������2O��1�&��h}&�@Vï�Y����jl�]��7CS�Jf���cO��=/"��l20J".�k���7��y�r��J<���w�]�����a]z��(���47����;���ᕜס�&��y �.��ɉ�W�,��yC(o��@t���6�eԉc�����-��޾A���Z]t�5��x������ p�\7>Bw��;gY�ecw,�o)����Եr�.�u�.���j�t�HLL�kb�T��ʻ��U޾E�z�4t�k�M��ԉ����>�iӪƴoJz�GL���A��חx8�1���u�ߥ�?�6m��]��[h� @�0�����jrj:�WՒط''b#1������ᇌ���8�M?�o�ҵ?�Q�ϻHž~U�M����ڜ�ݨ^���Z������a!e[�IM3o}�/�J��=�p�ej=��0�L����&����^CW]��?�Am��
�o�ZO<��<}(�;;[MA<��Nî��i�قo�g>��[>���];�U�m���oR�e�k!ѥ�{�)R?w965p��z�ޫ�.�\�_{�z݆��C��觲q���g4w�/Wԋݷ��t�J���?�JA���~�zW��-�i5wn�n�:;E�u� #sV^�i��,��S��*���`_�ڛu�o���}I�y�[Լ`=�2���1���K�#��5��^y�:'&�Z\�����n+G������}�z.ڠ��Ê�'o��Ǽ�jtL]?�^|��_}�V]�];?�SZ�ў�i���Y4�
A��2[��(��Q8Ú��5dk���zӟ~\�Mc��Se�F���-�}��VSQw���X"O.���>B�B������~G�3�Լ�;j-̆�/l@]Ѥ
��q@�~��y�)$�!tr���n��?��J�~`R��-Hy!��I$y�����O%aK����_�G>�EE���v!��ꭼZO?��Ӈ4��f�)��u��F��Z���Z�e��|X+Sy�����1�?����b]p��*=���}8�#}L�ބ���f��n�t�%�'�������S�gaY{֔�ӻ�y�zؖ ��T5'���$ej�՛�U��A�?p���{��D�f0��Cg�?z$��^z�-�Uڽ_�=/h��G5���u�;߄uV�E5����TN�,j,��M��Π�6,��ʽ��أ�k���7hq~J���g����O=��=�=�	1F:祉�/%�3(9��g20�Y$�>h[����]Ps�$$��G����V=�[�������N�����6�I�
����[����`�Qk�z=�K ��J�������%ؑ��jۏ|P�,��z6&O����K}�S�i�q/���W��U���8���A�����uK�*�ƕ�O���E��\]C��~ꔆ���94��;u�\����G���_Q�:6X����^}�Mz�g���ob��K����]ٴV�x�V�`	�X�o��_����������s�3�mȺ|&x'-{�K�U�xt<.]?��k��%�T!:���̙��gf���<���i-9g����_8�r����Q��|���W����)m���DP_?u\��>��Wi�G\=k�*�ʪ{�_S�^Է~�c��w���D�n�S��uM�iC�z�ٔ�A��ɤ-���MW^����[�a�PpWiB��ݭ�� ���t�ȑq}��t��aM<�"އM����0�\��� �j� ~Bk�]J�J�.���:_�YW~�g��i�yk�c��"��!Q/�ᇟ���Z�S�=6���-�B�<�'����^�+��-7k�UW*��T��u�]�j���ݏd�i�}����{���~ b�K�5=�=w�6� wUG{��?�����=�h�oך�68B�#�Z��eo�C�����ܪA�Y��ܩ>2ʗ�^w���N�� �[ְ{�l�ɤ�=��>��˳���\����f�ڸaT�` 4^��0������^��jg�����/��{���Kǎ���o�]�_�'�30w��So�cu��{���}�k_� t���g*U��.���ܽӬ��}�W��Ѫ7`O-5���Ƃ.!}JR��<W��}��I׼�5�?=���<�S���Iw�pJ����CO���������χ�	fP�t�I�[���ڣ���ꟿ��!� ,���7-��n�T����3/��K/P�hQË�:VK,o/KZ׆�5���n��;0�&�Mp��4�J*hk���举��1�^r����{��5ԻJS_��ک���:d#U#���1������ �ƙ�m]���M�ih�=���:zp�K���w�S�>�O��+�N��yUK��#a���+�p�U�����Z��%5p���vj����ZU�xf�^ܻW��I�Xs���Wt�Ϋu���kYX}=y.�T��7�g�*%6��T�Z;sFä�=�K]=����{�6�a��7�Wd�!�H���.!���r��������c��|Q���U�t[i<:����m>����RU/ �&j>�(�'s��:��G4��V^��������j���:˵�o��ή˵j�ZdQTfŘ��{���j���P�[o�]�G)?4���ЛSdt�l+��;�Ա�%}���YOc��������ұjC��u�a�I�R5�f��= r7�ݑ�R׾tH�>�O:v�n��O�g�j��-*��~��ЕcVo7�f�.��� +B��,2�'�X��+.�ym� ����ojziAS��f
�h���\]��W_���W��'T��5Wh�[��+wxJh�H�Wql0�	���}�>���>��>����#3ݠ�̂.��U:�O��Тm��p��X���`����w%vޅ�*�#{o4 '��Җ�ܥ��)�}D�cM�g^��C�����*�N�1;���?�o���虿���\B��&G����\m �A�2�l0�$��{�$�����R�Z�4_�i��>��rKe�U��Ѷ��֚�+��Խ����W� R�7�dU��4����~�6l�"���������#kٲ��r���$��iM���|߇����^/��	{l�,��Lf2&o��h�S	��IG����U���n$Xt���5��܌�1A
ȵ_������K�{��=�m(�<��w�V��ގ�
) V�:��QG�ޯ��w��̤ �a��V��L���4@���݀Uѩc���!�)щv�߆P�y������O��z�Nj���\ѯ��CJ?_/�^P)��b����S��NM
RL��cn�W��;��׾A�cҋ/(7?N
�V��}��G�kvҞѪ�(u̪q�f)j]R�L��h��YO�&t� �0�!M��8�koF�~���}��g&t�`�a#i�COq�'2<��vz�K���b�8�1^kk>��PeQ�u+�4��[�AR�v�V7�8��qO^��yH�ն�t�5Wj��W&�NS�h����N�aZ�u��I)����DfM������Ȓ�ȧ1�����r��ސ���0k�T�t��c��?�b�K�SK8�*�Mq�$��x�y��J<���Va����x5Rg�KS�N���G��,�W]��S'T���R򳢐������A�I"3?��o?��2���,YU�/��|D�}�;ܴV��l���: !hǓ���f��ׯ}�>��5>���6�*��|F��鼭������b�t������=������ݐ%����9�Z��Α�����oݭ��va�y2�~���� N���л�z��S�� ���9�L>��!��T7������N��ߪ	�"5^!��<^����Ҹ@�@�O��mm����}V�d�d�.s Tn�:=���:��C�Gg�v�N|�������3���PW�S���:�̃�m���sx�u]d�^���-�>�<uXխZ���J�_�|�@6��v�J�Ї~��4Xj���gsmƭ���џ|�3:����G�!�
N$�m���=�>���3::>�{��U�*�X[ԙ&a[�&M�2�6�����`	��	>�o�L�-kW��5}F�b���M:�{u폼��\���O�S	ֳE�F�뮷�k����'�� NHe�S�yM�}I�.�B����ʓ����l��t�U�rj	Z������n{�AE'f՚��t<�*��ï�R��֔��ⴥ�O��٨�aR���psN#�G��ǟ�酢�<��j�Mm�v���>)3��;4�-lq�V���.��������W�_�EU'N�>U4E,2 ��j�
0`���={P)���Ը&�w���<
'Zs*N�tN���7C��j�`K��,�����X�ϺI-�.�����]��Gt��E�q�Һ����k/W�W�o?�׿�-:�G�Eg����bQ��dR����iOy���a�%�ղJ >f�~�C�2���Ž�w?��ۥvH���ӟt������c�ҽ?�����q�P+���IP��"Z5���t���y��ۡO�xB�0<���z��F��-N�7������2Z��K�SdK^��W��l
]��[R5���0c z_�n��1{�׺;�F1���8,�h�+�Q?�'F&�3o5�=ї�5�D	�cOtE�:N�Fw ���oߪ��1����Ӈ��S/��4�q�ݭIX�G��ƂSO24���$��v�z�� /pY6R��HR��Y���^����ٗm�]�q���V9K����DU��݌%m"흃�(T`�U�c���ZP�*�=�*6�vx��q�f=wpR��ѤDPi��)��gK��06�Ns*���a�< �~�5ԥ+������hJ7ʏ�k��{��9 a�Y��6���cb�f���+��Tjg��n�id�V�`��ʙ"���2Yʬ���RM�o&�ŹӪ��N@:�V�L����O�`9����؇����Y"�w-@���pD�(��M�R�Y%�3�� F-�f�-K��Y*�C�<�7 wto�K+ZZ�.�ޞ���=�U5H!D��o9Sh��C�]n�-4�¤����
`�W�zź��'�yf�ǲ<��ܼv�m�cK�XG$�M���Xe�3J���5WPs��b����!~;6������j���Tk��CR�q��艮nE�FO��1�����f�5�lz���v�k5Y��c�#'�8D�,ـ��^�b�s6�m��٬���y�w�ށr��%��߯u�=@?��5���E�[�!�x �5d��^{�Y��2�}����
�{������뿬�����i?����H�<y�Oi�J+^���L�F�Uoy+0ΣD��h�p�Q���μl����<}�B��SÏ�<�ޫ�j���'��PwC�]ӥ�q��P\�.�";���7T��r=سR�ϿPO��]��!��D���O�N��r�+��eOO � ��D�8�Y����p�}>�$�� ZC�������{҄T��z"��p�2\�HZEuh���yګ_+�~��I����Sm�o���a#߂᷈b��I&M�{��4�X1��f��nyz�q���\�$�	���[�zV��y�	��jg]$1H���j��=+&�?�=<L��^0wgzU�(e=ʎ�5�Д.v "���o�lTOmܦ���U/<�i8�����N��*�UIԵj���ęidV�8�U��s[.������I��l;~�P��d�}<�A�����V?��n6M�£�p^��҈��bO���/��� ��-/p�|������]@�)�ItAπ��O��y.vM�l��	Iu��4�M�����sW��g`�a��2�+�I�5;0xM�F�H��	��|Δk�g�+���c0��n�S���Z�͒5y xinA�]�I#Kj?�z�0�m�A��s�7��o�0bg��D�_KK#ԍP��
�_��A�N��������O�Ƿ��Ҁ���l�s���0�/I�2��T)ꡁA=Z.��o�`'�]��yw�@� [ �����[Ѫ��~�����9�sdl���r�X&���A���I��ʤ�aJ��^ϲ��h���q0�J�#�浀�A[<[�����.=Ni��{�N��4�ؽ�@����WrF?qe[�&����g&9�A�Ķ�->��O�b===�x5E����Ԝf�����j�X���LЋ�Cэ�S2b������{�Rz�kB������:�P<P�ie��dk�)�0�	�d-�`�AH�t31*E#�H)�q8�����gH��p��V`g���m
����R�̟�?=;����: ��ӱ�iM�P�V�� 8"`�ͅ��p���s�1��nE�	�+M���s�F�jyoD� d�E�PBRY�ʡ�$J 	�5y(j�;�����S�`��O�t�r��q9<�x~w�����������ǟӆ���6��Oi�'>��w��x��	��ڴ�hh^�0� )|�$�r@����TC����I,1W������yEa�����5���� E�&�کڲ��aN�������N?V��
��1:��̽���k��tv�$�s:M�>����������v��gg�Z�)e��%85?�|%~��T�菫�y:������۳o� /��	�2[�,��\`'h(�&���mȅ��<_����ю�8��jqV�u�_H /�IRB��8�"ȏs_�u�/Ⱥ�@�OЊE rt�)n�JKU���]o����_�]W!{g8w�m��F����ЕW���L6�S���Y^���#H�W E�T��Wp��CI���S���upt���r��Q�_x�V�Ŀ�����z8ۣ���*]|���[����\/����=M0�'����[�8�h��
�p9�Y-���@�)?"����&�{&��Og �&�Vo�����U�K'�-�1&Gp��[�s�@�~�x&��D�A^�ЫN��'AZ��-�J 3\���6-���ح�=0̜#�/	�:�I��$���ey�*��$�zJ�(@z✛���4%ԗ��m��>NV���AP��u�5@ρd �0I���{��k��w�����^�ׂD�ȅ&��S�EgFM�L��� �{v�6��@w)��S:�P�~즛 �#�t�&$�2��9S�L�?���s�=R���۔a���t<e4��{��e�Na��~�;������Fx��K��4ֱM�������tp*���3�$0e��s���X3�0T��JeY�ߖ�a�8F
J���$��.�m~����Z]q������Q�y-O�J���~�#z�m��_s�2K�;�� ¥^B���G{���:cˇ5wJU�x-8��<��S��E-��2Я�W ��uz���BE>��`���]s����j�X�<l��x%玲�,�bc�S����K��F��x��
����<=� ���+ux��3-��a������YQ8 Y@��Z6(����C�1�-���c{�Wnza�μwG���j0n.��ϭs��En�Km�6��g��X�i(���zR4̵�_9�����������O�Ѝ���-�jR�z1K�Moҧ���:2~PW��M*=�$��B��.-w������.�0�$of���{�d�ɱ�41��*[��c�\��f�h���O�r7�\3���n��{�i��@��í��h��W]�i}��F��]9�xN���M����r�.z�T=6���*T�L���0�FjagW/<t�L�+W�v����켴�u��;�M��x��N<J���mݤ�[7��g���'O �ipdD�<x�6��PEO����O���,c ����(��`�]�w��= ��� v(ߥ���,3N��>�	���T��S��oxE誋��C��x�q�� ����?k����]�~���zӫ`��6�֎W]�x�ze�F���+;M�K9��i�}�}�~�^���>Fю�xm���}WB��fU@�g�!٠g�c>=���J�q��)�^��MBG�	�A3 w/x懴�4���~�ɴ����+r�z2Ģ*yU��_OR}w�J��+�89r9Kv�� ���L��}˳Ϭw�&�)�Y�JW�w��'%�6��e���2E�p��?{��g�5<ل������}�{�臄ةν�7#(�{A�G�#���6�0�����PŧIQs8V���S��ӰSL�7GzK%{p�^@�A����n�d�����O�z�}��^��)M���s�[,�ޝ��@<��}�ۏi������=tF�0wO��7?�����{r�^����Tc��������b_$�����~�{Թt�:k�+vf�RU*C�l����o?�ˌm&��`�/�ep
N��~����a���j������D͉g秴bd@�zT'���.���=�n����Jh�RE'I��k�؉�_���nPb�<�"�� ��P����ouE�V~���]q��gT��|WRcwݨ��߬��iRI�L�޻i�z��S���l^~����ء��g��0D�C��q��n�;߮���:o���vh��vv���Kd[�W\���J�خ��C�c��A����ؓS����ރڰ��n?O��<;�)�h�t�E �s�{ujF�KfC�k$qP�[����jL@�v�֌�St�l.�����K[�k!�U��K���[�'_��z��ө���/���bV���_�O=Ot�p}Y�2�*�t�������z���U�D���"�?��K���� ��!�J�[�*P;�ٽ��W�{us ��ݠ������!3�(A�P+�ך�ށ�U�����ӧO�/�։�/�A�+�n���^�C6�cnڭG.d|�� �՟���M~��6@hYNC"&��m;C}[Y�%��i ���W�Rb�fi�J�G�Ԃ`u֎)��<�W�uh���"�q�^�����ow�: ��f����߼M[��6]���J��I->�֞� �d铛�����/5t�ͯW���h/�<<�̍�ESr;��:K�9L��E� 5l]��\��>N�j� 4ؔ͚��m��jM��ڃL�[G�������D���ڟ* �@V���~L��7������R�L���7��&�mު��v�$V'{�fWD�z	"gy8��D��{w��w�U��m�u�kճ���I8��v�Lr̠�=����<����D�x8�'�({׻���w������*����a��?i�� ����y��~-<Ƒ���N�S�n��DpD%��M������K�=�4ʱ�B����|F̪��`f����^��#��a(�7��+ Y
�]3��i/�?�����~P�����;|��0�[�`���ZV��Sz��ֺ+.O%j=���ڋg�Rp��*z#�U ���qW��}�fnn�ٽw�넦oߪj�_鮄jKZ�ZR����y���7I�.�=n%�]�pD?����՗�ljT�~���-�V�Hk��"���i��a�]�f_���Ꮀ7���a�Q���w�R+6�$��lF0��)5q��N����;����y���oQ����,�m,r��z�;^��
@8pjB��!0&I�xx�TS������ʞ9��WN:��$�cr��
�|�u�+��^->�$:'3�ƀ��qtw��,&�M��TY�I��~N�:��O�h�oS��iM���e�p�҉AR� ��*=� 3! ��|NC�����	�R��ӕ�\�o=��q��о���]�^��8����z��~�m����~�l�K�,	p��a�$w@ʶl���&I�=�q9���9����`E|wVk��zgUf@|��ޤ̪�:�'���)���U#�Z��hkOF;W�\����/h뺭ھ�Z�����Z��Ds��4��+���$����b��,u�Af���5�S� ˘j����h1�Ӆx��ow韟٧�oz�r;w�O�q����.ۥ�Ks�v�R& 1������e��l���U�u���:�q���O�N�֔������s������������.�L��v���v!R��7� -���3�a�[rdC �x�g�6 {������N$�]R#�h�3�Mk�SyӰf�@�Ɣ[�V=�C���`7���$X��^��<�g^tӭ�̚^z�q ���~j�������G�Lq�r{�(Kbه�:� �66[�	~s����`x�q�2X����_Lx�%��n>z�x{�r��?RË�]���~<m���Rz��G]Hx���I�O>�&�ة��ƽg�Y׵��U�蹨�\A�E@���kMy�eTx�y/a5R��s�V�QE*Y�,�5/`hEދ+��-�}��G4��ER*?K�	�t�lܬ�P\W�p���\����	���Ǳ��λ�bm�ߥ��q���T�S͍��Żlj��F�G�m�EJNN��������OJ��VHӭs���[�2�c�����w�Ejk�����̹��Y�v�4_��c���|�6ʺ��K�rI���?
�h;�F�TX����,�y��ň�#g��k��-����Zy�0W}��gaGA*�z�vޛt� �{�_�=#�8��Sכ^���JM<̚,��Б����2���}�:���������r���k�s��";�s7Gzn��Mk�����G�n�a'��l
{�*�?���h��C�jP�P���9������������~�b�ޤO�{���˿�����@�{N���?�>���UW�����.�N<˩Fo��W���\���W��;Z\jk~������r睚޷G�u��6�h���|���a��ZڽO:�*�\d|���"`5r)-vR��x�ʷߦO�xBՍ�4�n����'�t�[_���'�#�y����g��1Q!�cd�0�]9�gK:��oi�XRnrB�}dx{^Pe�!uU��}��yQ�e�,�����}�H��`�ޜ� �A=��]]�����>�'6t���a˽�4�gg�F���Z]���ѱ�Y����uG�U�Q׎˶����FVn�����P�n�-�}z��Q��y8Z/i�@��<���Y2jo�0�/�u��	���'�d�)�8rYe�j0��/}[Qd_O��$~lve�[� ��`�7�3u��y�}��I�O��ĵ Q�,�l��oE@y��o�
���_��^��Ϫ�Ϣ�1d7��Y�ȩY[R�����"�8�Ԑ��jkn��� �+'4>I��[�.؇Y�W�;mOe�Wɣ ����X���!�����nZ�{�Ф�=O]Կ� ��<5��
�G]@��ڃ6�ޮnp1�\�^���':V�U͠_�cl �1���<��{E�>{�r�~6��ˇ���T�I%���m���jۛ(�(�h���xG_�x!���Šp\O�r�_�PP�����lIů~W����	���=�;Cݓss�8_�%����>��CO���,;�A����h�N�R����������'?� ���� �S�6�JLT���G0�9P�N6����p+$L���ܕ`Axz�ൻ �n�kl�z���O2�33k'g�~f�R����߮�|b\�viQ񬕊џ91�5�o�eo�S#+F4�7���y���u=)e>��Z�r���gu�C���ڿ� �n͗�T��'ѣ���Q�P�6�l��=!Xz�9�mD�^w��}��Z��h���]�9�,'����0Ӟ��T^�Z��)���J+�]��G��C�L
��z�zn��;>�^���_T�U?�GE�GC�,�g�2T/��2���{aU(��=[dv��N�����;��/aU55�I}灇t��7��'�����{t����٣�WD�3����54�k����Q=������;���>�͏i].�Ç�i@?�k�83���{)c�e�#�=��f	�d@(�S'����^����Y�����7�{�~����~n�n��.}�k���������r�V�f�_�a���rz�T�zw��-�Q2��?��u�qR�$��Yp+v�l�����-E6��K"�ʹ���1������@��y`��\=���L�8!r=�h�e��gU�i|���RC���6;�MO�俩�_�n�J3ϼ�n��cǕ#`{`=ͽB�?�4d���c���{K���+Ե0�.��U�,ۓ4��{?���~U~\��I�<ݱ��U�#�tisI� Er�^�s��|���]�*��h��ڼĽg��R���X�4�%�f�A-.>�{����26_�h&��Okŏ�Z�}�[j�!
/�����iizfRg�!���=uRG�U�w�՚�y�	xFy�0c}�&��6�i_�u��2�AM��-\L&�A�^i��$�V��<Y�YixR��Cp&+��R��I��k�A�%�^��魊O�/���?B"%�:���=:�Q�4,A��H��G=7ڠfVB�����7h��VNQ]��M����&���V����zj��J��Qַ���\9<U�v������ {��F�u~�F\B@�BJ���7C-ܭ�P.� �!�Wa���z��!R� Ɩ�7i� r���jj__@00kcF���كSضg� s]���-�#�\�y��[n/�le"N��3X�wݮ���H� ; ߨ�~�
Ƙ�����+]ҝ�޾a}�dY�a��5�Kz��s�<�1��t�����4��.sGo�]����j=���#,K S�9��$��R�Չ�6\�Cc7ܠ؉�����aHIRww! f�dx�[�,�=���x�eg��G����7�4}J��1��+�B�	����Aw���r��5:>=��X���-�� ����^�3����� ��SP���&mz�O��3(�����?��W^	9H�ؑ#*�����|@�}�꼫�W�s_Tc񰒅�*�����Ef��u�A-��e�A�6�$��	���G�v���ѴF �����M�<�΃�v�Ҧ�J��okņ�������+����G����-;xT=dU��˿�����އ�SaaV�}_*a[��-��zl��d��@f�~�!p����ŀ~ȣ�@"E�c�в�%�um��߄�a~�|��&U�zO�zMnP�mد6Vm�� �|��z�s�Pϖ�Y���!{�N�~�M�N`Y*k��v��N��?+?�m�(����O@m=�©���]yM@�ġ��'i@,��	�B�<���^�Ә�M�7}oꛂŦ)�X[�F�H1�����۶<���q�y�&�]y�C�6zP})N6�J�_z����ʬ���gNk��g���Υ�8������Ɔ�ߝ�4O}
�3����Z;B�s�F֌��g>�m{�SgtH��-`�L����;��/'kUl�������J�=@��M^��.�
�����	��,�S�B�b�T��������n��_� ����'�F����Z��+R�\0�$a�Vi@(���f������p��aE%7�!�8��!���޲M�gt�/�K��z}�_>���NX��7���lӞ?�%��ZSS8xF�j3�����h�sQD�EXv�9��	p�h�~IG�w%���ؒ]���MiQ��Vm`�s_�bHc��0��6.�U⮆:lb��Fj��3��SA�.ى�>�f�[�}"�|�3񞬞҅�ⴡU��==/˒n^3�W�~����rD�����\��8{H�2J�o�9�-��J�ʚ�%�Q���
H#[��2��0�\wN�4�\���� |"g�sx=�!�'����7m�����}���Ij�'��9���q7�"F9��r�l�K����y@��]wa�6��8rv���!x)�?r���$��;���/�7Y���.�@*R'��*�����j�-��_���~C��slYG`n�4rsM &Q�T�YQu|��'<��IM�.�;�M4S��	x�pF?����Zv�q�����b�z=�տҪ빧�-n}$<إ�7�׾�N=�7���ko�����8�A ;t��k?Wl�X-�S:���ˍHp�`�Um@W^z�	(�G�=��,�sŽ�$�@���i�-M&�.#����!0a��J0�����F��z0׋X���$��~ʜ�6��(�2����W����i�퇠�v��n'<�h`
�A���xu�J8�r�>Ҵ�O�J؟l-�c�O`���圬�_���AO��x�;R"��R�3�N�g�q����
�wE���E�%2�����dT�f�|�P��d=����$�{:p��������.X���fP*JU�-JawՌ:	H�����e0cOc��3~�vS�غJ��T��xK�M�ng�!���(��w���]���~T�RI�)�d�˨�o��V��AV/�^|�}N��_��'�UU�0�k��TdvW^�D@����)3����ϥ���-;�~'�>�C�* ��Q��W%����[����3%����<��u?���.�����o�E�o<���gH�1�)��<hT����V���o�}J�j	@�����:�� � �D�v9o�к�*M=�l� Z ���`��><W�{�xAYkl�΢�رM$+:?�UvnR+�J���ά&j���A"NŽ���6VwsىHO���NZ�� �
�ݸ-��H�:� �<�ғ%u�g5G��H�B(����e3��'�'��lf8�]�n/?̃X���c��xֈwBD�H�À�@� g���*ׂ�F�R?a+[*���+������8��x��-�5fSm��.a���3��9!#Sk�X��vg������W��ǧ*�����~ģ����qV�F�	Q� h����s�mH�5a����c1���o�����͜�$g�%RU��թ	�I�y�3�&(���s(�Pf��iu�m;O��r戆V�>�����ji?�#�B>�����Z��N�߽?�O�& A[2�����|!=�:N����v�M�4�����s����M�b��K���{�Ӏ��_�َ�^����wMY�։���:��gEA3�����<A"ml�cw	�d� o��#0Kȑ�j�2�w�P�P^X�ǽܝ�7,�6��ň8�=�L
�e������V۽��x�HX��mE�i1Q��!��˵��K�{yf�T=�+[���|�~A-��2���Q=S��[�Ы���u�#sK֔�>���n0������� 吁��Ӟ]UŞ<�,��w�����锁t��9����c]�'�7��1�_�`���pM���������wCu�8�}5�z[I��ΪE��ƃ^O/���gՁ���ӟi�{ބ��kߛ���.�}Z�G��Vd��S{l��;I	*D��{B�<��4�\�T�ԃ_��(����t;�G����'tt��Z<5����K*��ŖpΞ��<�[Zӫu���;�K���:�-�c���4�n�"[����%��*�/�q��v,�G2�p��/E��x��z��Z�I��gx�l��J�#�8���pb��֭�Y��̪ؓ�v�k�����ʘ@ @�9ni�s:��$v>�Q&E`�"\���2�!�@��Dq!~���o��D��w�bZ��\o�	7�6�����f�J�O:u�i����36��0�fܺ�~;sxX2u�Cz�� ��36/83�s�wSN�ρ��YM`���HVp�"������ �I{%��{a� �a���Ri�+��X.fS~P�Y��{%�V:e�&��q/oڔ��{��gӄ��g��50�BW���G����~t�,u�u˼�/����Y>�'"w;�91I�s�nMO)>;�>Eb���줚ӳZufJk��U<yZ�R��%-<�_��l3Zˠ�~�dk����'(�h% ��B��[|B�)�^�հtPF~tc��u�tW�z��cO�SP�t��E @�H?�c�&���!�l�;��x�����
|��]�wv��@m����Í8�@��.�[���=O�z���9�f� ��6Fi|�AK����0 ��{śm{\���y=I��G[��o��O����:�_}��Z�O:��w�I�n��6U[vSU��g���
��?���K�~l�������ae� ̚xV��>7��}�Ti�
��Ud% �㝀��0~d�:�a�+��Do8��r���:J����R2Jr4�١�{R<�Eۗ(��fH�tF�k.��廴8�E��AwZ��oH��SJ_�K�K/s�}��
�� ��O���3j�H�A�Ъ�j��0�&�6��	Տ�Q�F:S,�/�=Ԇ����^|� [��_��R�'T85��\AERp���M-9��ǞT����~�9��3G�C��2�_����ȇ��٤����i۵�����4��s�K�߾�y@��L�EF#���B��b��޻�T�{L/-MiǍ�hsyJ��gՋ9��#->���u��wܦ��E���Vn�R=OT��Қ."�� �-]�\����c�u�N���*2��	~�E���j@h5�?7rl=�.�i#��`��|�k9�����D�8��K|��8�Z��@Z�k�k(s%�������c�{M;�1�(׬D��d�� -�V�mo�҆yt�U @���� `[vL�	~o��y��zqp	:�o�e�Xl״)�' V���t����-)X��s��g�a��S���"d.�o���/��V���x7A���0��?���Ĺ����Zx���@x6�������~�}9��q���=lo�q3����m8�u���'��cJț�Aɐ]yk���6��1�d��=gza��﵌�ޒ$�i[2�Y���urP�eM	�5��-Q�Y2�*�
]!.��ߑ��;�;<���	wQ�4J�;6���s{=]_�L�82r}�y�f�=,�v��f�l(?�������-tIp�I����Q�o�ے8����F(ڟ.�k��O�3�_B 8�NV���e��@���U������.��[���/*@hƮ�R_��a�|�[�/=���z����{����sf��������D�k�,���ޣ[+��Q�E���Kꙛ�� �T��'K5�K���0�?Snk7�$�a�q2��0�)��p���FDӵ��!���X�8r���@�a�^H9)+��l�6Vضy["n��o��>����l�d�V�zUuW�_�f�`ׁ0e�l�OMϫ��ru]}�+:��.�2��]%ލa�q>@�ݧ�u��Sϩ����η�����j�
۩�ϰA �B�?Q���+���"�u�r�3u�� Őь9%��1�tw`��2��.����o��}�]�(K����+oy�VO�⿓W�4��N!�30$O=;/%=�L��=���|R�GX����>����Y, FӉ�|�E-��|כ���>���1�.��-d=[`dM��W���[2l#�H������$)�g��З�i���.3�p��g�H������I�4�.�d�w������N�Å�#�w�e���$�m?���خ�S�U��3r�Q���N��-��{u�;��]꾇?C��z�	� ��ӎD*Vq����vw��d���7�9p:��f�7G.�N�+�+F��^�-�P�I���S�U�g(K�K�#���D����=tNB�)�7����q�)���$�ɼ���z�:N�"*O�m܇���6����8�\]�ɑ�r�Et?�N8e�md�o I��wi
}�A�~��׷ě�0�dSWNs�����)ځ�{��) �ȧ�rTAn� ��[�2v�6���&�r;h+����p7���x'�XV���9����R��:�<۴����P��rp��z�W�˜�������~�@��w.��lA��ľ��uL�à}o?��7Z�~����%�z�����>�H�/���h���4�z�����}\?�c�Qp/�k�e�_����|�U��Ă�;7)��%.�o?���:l�U�x� 6W��<����w*�U����c�&��b���HR?��>���ϕ���U����PM��%�;�F�o�����0�y��z�i�R�=�7苑����(�~��;��׼�̷	a�CH ��������ݧ̍?��_���/�^|?��������� EY�֩�K��5�Ά���M�k���/<���)i��c%�V@!l�*��;����!�"�!�9V�j	�.rv����h��X�,҄�EQ���D2*F�0ö
ɴ?���l٢�:�s�Q��)j�F�2I��Bˏ��h��D��c������ܧ�58]WV��[��"-�aO�F�d^V���*��xvV=�:����Q �+.S�����\;D�#T�zF��
���e�<�H_1\�i�C9����W���k�� C���,
��'����`��|(<�q�3��׍�� 䁩)X�o��q3�͐��ݕ���������P��\���vp��b�=�n�W8�o\G��R�y�̩��<�3���z��FWZ����S���{�Dt!�K�ۇm4Sˁы��Y8�����Mq���0O��+���gp�PgW�A���z�q�fM�?�纹���u]���0�km��1ҧa����+�3}^���" ��.B���'�Y���e��l���.���i{���ߡ?��T1��3[/�������0�W �U��^� -"�$Y��S�"�����'�Da��2��к��rW��� g�3�\��ȷeY�Vi3������=x����>���,C_���݆L���8t��/��/��4���H�
d���������G����^�h�܇�gw@6�H�7���*�7�����id@��b�^�ٰV )7^��x���;ީ��C�f��qu*�gJ)u���u��q��[�k����O�,`^kGf੉ZR��������ǕڰF�W�� �`��1r�0n�w#�,3T���e},[�9-/o����S+7 ��Ma/�V�k��)�&�(u�nE��)����R�9��z�K�m�ǞP}�����5�Z�� �{�Qs�Z�E�`WR���"u��!XQV�����& �(	�"��iH�tp~��u��'��=8wg%=�I�0B��a< ��=�fbZ{����,"�L4�G��XM���[�m��J��&�X!�̤ts��5��F�����=Ktu�_�I��:z攺���y�m[*k �$��"?o�8`�-�S	u����%d�H�x#�Ч�vK�b�c���a�h�S��"Z�9�>�~Y_�yߞ>�;����|p���Y��N^F�U��p}G�*�x��ۃ|G�YMFaZ�z�bM���*�o� �â������_�E�lt�BX�!�h7���t�e���3��̆ W?���l#�!�6���gĘ����y�t� ��3AX�s-z�+�X�[�¢�o���g�l�A}=��`�T��9JX��g �����/����=�!�;8�ӿ�<#����/v?�q���<��ߙ炅��� =���T�rͪ��ݺ��%�5�h�����)>��&��x
?,���͙�~[Ǒ���m3@z�JXXc�������t4�ҁFyp�f�zwK��xv��r񧷓^��@��o�|�����sFh��
d5�c�ii�[A�$K�m�L�b��g��ǖI��i��!ξj;Z�֢^p����o�������z_�H;�{s>�1
�V;�:��]�kM$��j����~���I����Vt�4���Z���'&4��*^��v�DXD�i�T_Pl	bZ\Ta�A���Mc�h7�Jj9v����?�W��-*�.*�nD���W��Jj�TR0./���;oS�P�`�K��>D@K����q�>�?�Y� �q߼'
��Y˶�~�L!y�GgQM|�཈ Sq��������{4\>��K�?[R���/P߫�~���{�`օ��Wm�s�#Ĥy�YE�`� |b���H�lC��d	M�0j��:�ʹ�Ѝ��1��w����0�0��b�ˣ�6���V4�A^l��%s̧�_���Ӹ�fL��f�4-���$�۵��5����N��x�Qid�xfV�j�*�P��k��ϛ�0���ʶ��/���
����k���fA�5���Z-�8��r+�7�zg���%�y	�Q�2)����b~�=����~����rXDR�D�v�Ct�F��(��k,K�se/Kb4��s1h��;�镀 aU����`yc	��1�,"���'VU�jY��ĐE�x��ڳBl&T��04����,�,�'��!:u����x��}~�MW��B?�gR�O�s7S��	 ��1��z��m{Z�U5[�q�݈a-����\�fb�e�b�z0�/q��{u�!�{ey1
�����upq���#��7����՝b��Cjh���=����`U��\<��U�Ml�Yj�������L�n�wc��N��n=�� �G4�<��{R���ũ�&�t=�4	��2�9 {I�A�r�F�ck������ �<o)l`�C!\M .Am)#�^��9�>C�Z�g[��vc��T�&,e��U���v³��{�j���v�)�H �l0���K�r������CK�=����aa�b����v6����g��A�$�h�{�����������2�ҪŢf���rf\��%pl^�����E���y�|x� ~H#��������]/��}���j<|�2�7k�:K 9H�
z��'���2�l��D�[6����/�ҟ��9e��OOlp�\(׾@�O�8�aB�S��^�I~���d�y�t�8赩�	I>���;�O�Sg��^Rm�1�m�@�7�&����+��9���V�D��MUR��W߆���V�QC�1S5O�¹�'_���O���U�a�r�<��L� P<[��&�Ω�0��/h��[�kM�f#�:1�Ў�_Z1��i�����~�w�4;�|� ��q�&���jU�퍺�5�ו�ߢ�����i�u�h<�e� �q����m�^��\"}*[��V�hZZf���ʤu�ۜQ0�}�,�c��lہ�$�9���D&�fڛ7���7(��6�ޠ�\��u�v8i
(���8��b����q\{���z_��.�����i��=�|�b�Èk�>O�@�p93Z�!P�нYU: #�P/�O��!�鶺K���:n��tC+۶Sŭ��0�%��I�ͩl�9�X�h(��A��-�\f}u����0��i���Ʃ�H�@U�u*"���m�[f�D*�E�<.�Yz�~K<�x��Y졘���[�����^�Q0HXMR���'�eD�?*��a�"ë��U��-W�
p4�:X)�C�3̖Su��<���u��H�J���^�s�%l� ��a�fh� ��0.5�N���,���w����&8�B&��nH^���S�q_�aߔ�L0���P&�s�خm"��������B�u?�?�m�e����}��E �>;G�f{�Z¾*�2�_�R.��neԗ���)���|��� S=�R��'��g�6W0b������[�3>�2�B�z[�Z�+l��n9���p�i��8<�3̵�]GWH�v^������˱|�F܄�p��DVǱ-g�CzS�Y��" XM�5t!Q��.+��[�{���7�����~�zM��>���}U+֯��+�k��.�Oi�3p߱��ѕ��1={�Z���>�tkQ��1:y&��"-�|���[�ɴ���F�&&e5Ef�tg���bI�
�:����)5&�'0�|��mS߭�����z��Q^���}>���Ύ-�7�e���Y*I�f�b��)�<U�L��9�#l/x�`�Zܗ�ֹ��i�����5�a�G���h��u��y=�/���Ǿ�$�5����tx�ٙo|Y��>�<���G5JV[��B`,�h&��b���O�[ٮ� eS�>�����T0������GfU}��o�"�DM������/=� �`y�;�E<�>\g0H%��G3��POSQ����L��d�PmIP{�����>߻B�=�?[�E�.j?�1�ADd��o�!Y�^V^��&��j,����:�a�sI�#��eFh+p��d$�({0�=���%;��%�5�ugr6b�a��lH}`�q��Ŷ�9u�I�K.�u4��+;Md�������� ����D:0�
|�oUnץ�>=�R�h�չ�1�_x&4���C ʇp��[�
��[��
9r;-�5yF�{#u=K���pWVG��7ܤc#�Y�R��7����(x��P����S��lE~h�S���
�^{����L����S��~~��?�_��E-Z&��b� �l��w*�~mXU�E���e��O<C6�>�$�㦼�بv]���Y��M�9�$,;S��gt���<��� !��}���Z�����9yJ٣g�����/����g׸+��6��57�k�VM.,�x�Z��^��U�O��z�Pf��{���ٹKk_�� ��"��W=����z�@E�xZ��=�*��ש��<d���A-�5�0���r�|���'>� #��ùǖ�+H$�fi�E �"��LO�=͸�Րφ3��4t��X6uw�f�\���d��y�d�xe������t��l�f�̃_	aj'�qnp�e�K�lc&�m�oH�^N�F�яo�&fu�lF{��2m�|���k2QL>���*F���hux�2"33`�ϭ,&�H9D��:
�;U,�pQ�2'xڱ�D�y��n��#�1����8v�q��v�ny�6�ɟ�=^y}o>l�|�}���C%�D�V@˃ �����Ql1�P5��	���� 
MO�w�&�~N;̄l�����*�F*�"(��r����r�ֽ��a5KJmڬ��N�IahH`�𪫕�����K��Rl�z+WH%�[ӺL&tS�Fx��������.���ԑ���3_���+�!��,���h�k�1���}��Ǖ��t���u�їt>�7�j�qN� (�$j��0��� ف.�tanب�Dgo'���:u]���<����������p��!���#o04�m���B4I C'�8N�� r�����Q��������1s%�L
����IZ1����ê��t
���W?�ѣs���hf�$�(��h�V��7+z�uz���C�� ���KU+�U9z(<��[bx�x��O?�^E ���>�RF����7*rbF��)���A����uë�8r�a��zJ�����0�����A�Н0'���Z�]�*~i�&Ƨ5�=�Y���7_�&�s�����d�6�{���'?���*�~�iM���.,i�ڭ�l]�^RG��0�_�W|�}J����A�g�Nj͎���cO�u�zU@#�jɼ�zm����%�97W
�5���Ҟƒ��� h�u,��'��a�+�gu��50�ޝڰBݫ���ӏ��a���TQ�GީJ:�S'N�Ey'&+w�*�^��O�$ξ�L�~^���*��[5>K &�Ⱦ[�I�u�jni^���jC {a�g�s� ٴA׬���h�����7�<��ħcO?���mȷ%��/�տ^��U��kǗ�b�h��i�����|�Ê`�I�hx�W��q���:���q �5�d*&U5l�l��il�O�Z>��m{�'<tjd8��10���'��ЇP���W@�h"�A0#�S��U-VT��H��/@x�?/�"O�l�����fM������7l�i�L�H��4�L2Gƙ'��脳v��+߽~Ŧ��.����#R\���2�G�/�A��f������u᜗_��zM��P�ྐ6P6Q�B_fy^e��g4�k��7ޤ�57�q����ڥ��W*��B5{{aH�J�t���}J�:a�(�� Fe ڻF�P����ߥ�q�?��Ξ>���P�����%��� o9[�H���O�cU�B�r�\i�5	�q�fQ��s��ϖ���u�����{-m��Ă�m��6�Ɇ�nZ��w]���i5J����G��4
9P8��*P�����h^�K/�ȝ��y����&%n�F��*B������(9�ޢ�2��bKU]��o�)�	�<כ(nf�̮ۣ��y�u����U�+v�j^v��ut�,,��u�N�܌k���ppw���
��My%b�D� r�]���>~/��&�*�k��h��1aF�U];��mo���kl`8<㴃��_t�&�i~��ޯ�C�J]~���b�pӽ�*W+��sj-�5�u[x$����3b������S�H�fa���~5� @���ն�.W��f�𑐁�ȸj�ƴ��oГ��"+��/ߥr*����_�Y�LV�����z��#}�v�/�\G�8�z��MY��[(k�7�V�k<Uӳ�=X��=?��N7vzHYP$���0��e���	u��3�6����j��ޡ��E���^^t �ё՚�%9������;�����w���){LY 7�< ��;4���RV+�*dp�o�Sg�yM�xR�<�D��L�*����'N*�s�Q���<�;������dJ�'ߣ��AU��@��֞���ư�	����5j���o�+寧������#�s��ԬO=�ɘ,gmǆ&Z�9~�s��O�w�ZCê���;ܥ���b�0Vp����Te�1IX�d�D__D,�@�%��A�;픾�z� ����h멥^*��Z�͛&.<��|�m��(/e�E&��8'`�e�v(=@� ����d�*���Ǟ8��^�Y���K�u���̒"x�~��v��p+��O��&M��咎�����]�z�[l�J�W	����f�j+G);��g3�O�����G�L`���6�I�o�}y�������+�}��~�B8���fNq,��ƕ*���J��59�"�WiF�$��0?C1�c�қv�ۉ/����b"�W�S(��č�g�͑�gq���Ϩ<uJ�E�L)2_Qf���N�U��AM����7�ė��tc��~1k�W�/Sn�O�n�Z�m��ܼ.۶	�V��=�Ϝٳ��Qv�i��A�����ў��*,�:�Z@`��[)���rP]�y����Fu�whT% D�y�GG�y��	��tJ���g��Lb�����*��\G;�Q�j���0�����:Ɠ��Fu�Ѓ;/W��M��|�w�����J^|��ãj�W���A#�>��A}�o5a/�J� b�(�w�	�i����'��A�~�M�g��{a��d���ʨ��/<0�0=��3Z�;��A㪿tL����[/��2�`���]��.�3/�Q�m�Z<;��s�!�HX?�;n��y�vH�������<A���p�U?���g�)�1u��ߨ�`&�?0��RE��ܱ�Z�q���$��)����jr�.�l~P�DG�Z�6����3�̎Ӗ�4>5���O�~x�
m�ֽ�͗a���d3e��^EoǝĦ6�Sy����p;gc���ui~V}�i�����g�hld�=�Q��Y�;��,b��nR�����-�����5���n�X����zp۳���ݽ�}z����;w�t�F�b�
H�l�q v�'�q��$�I,cف�!ŀ�c!$1H��`4s��;w��^N����{��Hd��s����_�+��~�|K��e�5 �MF ��~P�
����wVU�i*�Do��O��_Q��㳕�Q%�|��<��������ԫU53>� �kהY_��	��@��0��&U����;j��s��Ȗ�:r�EM���O�|<��S���{I����ib�Ο�����/��g�@S��7�I���<?�j�<ÿ�K�vT�~ɩ����N_�=OA�Ɩ]�y{-�t�d�e|�˙�]zσ����A��R���␉�x��G���o���������=g �#�}�Q}��W�ި(6�Pb|HWj��I�U�[ǫ��j�=d��r��'`��y��V���+�n��x�(�$c���������^u��2�=w�GO�|��J'N�9�W�\Ql�|Tk;dl�82$+�]����'m�uտ���7����4�K뒀S�����g=q\'�~4����z.WP�!��d�(Zᘯ��MR�M�On�vaK�TC��o���GU�`+���,)�^��,�p_���(h/�6A�����@����c�`y>"̰n�8����F�5 ��� x�o��E<q��J .ё�@�m���_�M��e�کiϋu�{�S������~$�A"�6���/�u�yM���O*34�sD	�߫36��0�C��N��}�
�$��5R=͍�vbz����� ������c��|���9��ك��d�N�S�|`�p�c ���u��W��;j46B����0�J?]{��m�en{�)�K!�TE7Ό�;mm�M=��jk�4rTB��z�[��{ަ2����R��W�6Eq���0����O)Z������h�{g�9{f;�c��
�c���m��ֶ�~�{,�V��9ovz��	홚3������]U�^^-i�=oU�(~��Á� ��֖�·Uc[�mu\	��V�͎@R�kzjF�'�k�C���8���c�EK���.�@��K����S7QЁ#�4>T$x�d*c����������{#!Nރ�ϼ�Q2����s\)��K���5q����s/���Ɠ0�N+���#*����%��:�ʖڵ���;���_[�/�[v朿�>�	�w�;���)�muʛ�� GV���j�f��w����%
�?t��������!-ş}N����J�sZ��͒	�g��ߦ6�n�\�hn�^5Kk�=q^]�pyc)�.�Y�WjyY� �ۚ˫�!�<�W�k-��o +g�w>;��~��Z�?��oR��o��W���h(8��i\�hL�E;�"����z㛱a�cӭ�5%�+j�G�����}���)����"����K��o "s)��!|��k�����:Ɂ.\|V��*���d!�uH�G>��Z__�ȹӚ�Y\+���/�
����+d�km��1Eh�������	�ϝ��x����G�"�����CPs雅3�,:t疚&�����82����{"b�����o5v�i$�Pm �؇a�9�?r�:D$/�aD�4(��*�+�,-kc{0&�ݣ�ޭ~,S��N(�u�4�i��Gd�D���(,ߵ�;D�L6�,Λ�=��4g�0��u�B�0������a`���4����<c_�{���ÇS��iV踁�:ݴBӄ-�������]82����N6�j~�ɏ��ZݴN�s�F�jdj.�����Vu���5<\$@6��8��c��~�[B���&��Rj�%�� 3	@�!B{qZ��h^�}oU��~p�Q�gT#�1�#%8,b�Uէy�'a�����軔�ɧ���i�`wH'F�H~GƖ��77�4�k���F;<������j �
έ�����*7���9�MM�n��د��MŶ�]k�DF���l���E�f3*��L�l��gJ�m<�p�悒�#l�r(��7ל�r����2�q����xaV�VO�?���^@�f<�V�}G������05������b�	�;Ue:�'lܬ�D ��0{M��ľ9�;� �Ք��2As�`��C>����W� n��Lڣ1ltzϘb��|l�;φq�$���1-��c�5��M���Ĺ	�]�Vwc+��l��.����>�Q�~�G3��?�,�@��Ӈ�x.��0N�����h*�Awi�F&�����*�V[��y���E��;�TR��E���!	��1������j0ro���!�G(�Ґ@g��#GT�C����c���w }��:K��B����!�����q�ҙO|P����]�7�(��D^w�2��wH������������*�񝄆���{���<b �r-2V�K������LT����}�T��_�O0o 0�=oR�`� X�fp��F��Y
��0��Vc�ݽ~�e�l�!�e�}(�Q��$i-xL�ΆZ�����Zƾ�Gk��K�[N���l.��/dW�?��J�M=x�-ʧ�U��<1��#c�'�v	i��[�]�G Q\>̝�po���3��ۏ��6�Ǿ3�jN[�	��wݭȃ�=��ݬ�V.�]�IGvvt����°+�-�}��Z_,Kˋ�n�ioH��]C���qM�P�i��63�,idK �Ǔ�S�_��㈦{Q�eF�c&�*��_|$(&<��u^�4���La�M����8�P�uGq���	𵜮�+x�h���]"���O.��g���g%f���bG�=�upH� X���l�Y.ig}EK7nkkcv������1��f텋C���mi �&�>߽A0j�D��C������1��2�g�m��V%�썥��nkceI�j	�m�ӻn5`d+;Jn����MSvw�z�/&��
�=�ښ���?o��&��F,\�R]lQB -ѷ���AU����iljX�I]�W�MST�ڡ�.��>��̡�r��*L=�.h��A�֢^�ܿ�ޣ�Px�z�-itB+�e�d<s��j��ϵ}�Y�a+���϶����L���Wְ����G��=�g~�ks{��������,޸����Va�u���<vσ�.����W�H�d;Q�OY�R}�T��s���h|j�ν����_h����d6�-�[ǐ���7ԛ{-V�]F7(�;sD�����ʂ��0��"h.wTY\P����!�3g��Gߧ����U�7���3 ������*�V�7�!�f���	;xA����ѳ�g�Chg Ug���.���c�&Y#Ú�3���}I��E�:��¢�8sW8N�Uoh��P���Y�%,[L=M�kcK�{��4���Z�g�}�j�`ʿJ���rD����O���XQͦ5���k�֊��������-7��:M	t��M�ц��IÍ��K �=O������?���{4�,��zR��8�D�=�"йq1�Ŋ��.�0�F8���zaL�����/I�[JHkzcEg�鳓E�33����B떖��Y��~��"�Ε�"��B�	�
����j�̚�z�]�T�Ȝ��j���!�k �V�J65��eF	&��~3���)M/^S�`v'C8��Q�|�'vOA�����+�h�_Q����HL�O|R���=p!F5�C��c��s�,��S����P&��chCڮl+��e����b0�.@�(]�o>�CJhvg�&"�g�C�[��A�h�`�)��0�C;���Q��y��c�.O�������M0���)��S���C��9Cڄr�`:�V�/���,�4�������jdr_hCq��sxL�����)�²Vn^U<��wj��Mup�)_����|q���đU[��:�����6�O�T��'�`��������&�����e� �n f��aU�w��(��+6&���gY^�)3[�砝Ռ��^��"/%]#~&7�@^Qo�@��6��"�s񲪷�*�%��{R7������#������q��dOן:��g.��ڋ�-(����W���}�L	6W!+�tw��ʯ\Wm��
����_�����1;:qp @�@{j�vC�������uj��^���K��a��v�Y3�(�A��K��IE��;�ũ6��n���9���yDb��P^m[&��tE��7���Ό����_����W;ZE�Y���,�x��ȥ�j\��^}K��G������ڹy1,�DhaIq�B�aH/i���b��k����N��^�6�  ���\��eC��ޝ;*��$c򆣯?������z(�~��ql`:��ȋ�!]m^�����;VT�,�֗��q��c/0�q dc@p�6~�}?q��\��}���d1�deS�W^�����#���~Y}��X{�߭���intHՋ� um��:�ةm��V��H�K��-��I٬ul2V6���s8�Y�nV���	���r�P[Q�T�[~�3���ջ�<�Å"a�>z��7@r�K��	_o��P�^�Q����}dxF���n~�;ڹ���u�����5��\ӱzIG��M|��ZM�qP�k{E�2�\�����E��k�Oh�C�U,5�s��M��X���o��k��6�t����A����Gu��� s.]
�և0����?��@*- h�����>�ÒH�Z�D������@G`c����Z���m�--�ZZ��%ݾ}M��;:�γ�;q��|�qE��w	{�?��`<6z"���AYN�2V6�6p��
4|wӊU `�;:��^���<�#HxG�k��^��
|!�R�xZ��n��s��
\��i�z�����ao��+��j;�������*ї��CVʳ��g��k;z�G?�Lj\)��M�O��\]�{}���V�����E�����ŧ�W�o�-��c�ڧ�i=h��4��сV���Ͷj�j���)�������5���aī2�J[����ݸ���_����M��3?+x]C���.��W��������ݧ'�����]�,'�ذk�#��!�;:(z�Țp��u^�v�z�	$I ��X��h����pt#mp�	yA��Lfi^5��$�hG��$	F �����rM�R��f@{��uhW��v�Y�գ��BS}���J85�FpK �W븺���듑�L�� ��Y���Aύ�)�"���RŤ�G�!��ϩ{.�3-�˥
�QdH��jJd��P��&�M�v�HPV�U�iA��X�`YěQ����Yz)!�*5W�&���K"��3h�܇�O�e�8)�گ��'dd���7Vz"A�=It���a�g�{r� S�Ӽ�C������k4L��������zlg����O���ŏ��4��?)�̸	\�CH]�KJx������J.|�^�\G�w#�O�Tu���P\�6�6���c�쳊��6::�!�/i�k�׿?���J�,�؆3�(5�`ʡ�Tr��,��e�h}m"��R)�o{�(�:��7�Ѵm'�t���2�	�����4F�ܫ����/�c<{Ǧ�g�܏(�c���h��K|���n7�	ط�;����p�	���mo��x��5�}���R��P*�U/�G���Jy���4��@��
��1 �s��Pp]%>�G�o�Nqj��R�|>0�!R��b�,��&f��52y�����ʶ"0�w%by>K �T�1%�d+\7�10�@O4z��F��Ժ�m�VJ+����M�� ���}/��#CL*>$Ļ�p.���HBg�)���v�xѰе�������T%����e�]�jp�i���KeB@���}k���&������c#��&=�O�܀���bfYpmҷ�;-����_������y����A$J i���P� ��e�J�H��O~��Liv�u���7˅�I�D����TK\$Sk8rl�ip�I�;�� ŁlJ�3	�OGu��O��I��X2K��gJ��9��=�1��rI=���n��,N�o0�g`u�����ni� �����u�w4W���l�t&���lu[���B��`���<�쬋�c؉�"\��O�Y1�R$�R=%�k8�}��ؓ���C��XA
����� �����t6j����&�Ϊ�z���3�t�Ap0Xys_V��-v��C���-g]mMa�' �ʓ����O�<E ;� Ǫ��G��ޓ�A}��^�R��^׆*��X*�!�f�td�� �"�<�>H�'!4}���ܮ_�)Rq ?���K���}�1��FΎ	iaC_�������KI��D�w%;� c���o�$O���W~����O�o�����җ�픲��fNB�δ��?�f��۵]�u	�Ң�f�������*zDٿ��J��!y��FO��U���fu�|����㼏��W���}{���.�>}
�	}2F�.��!�䗯7��R
_�b�k�5tn�9���ShB���g�0׎�*��C�L����!,�k<�L�)�-�2�4���d�w?��P��O�klvV׮^V�Z��̴���bS�d�����"�޿�ؽ_�O3?�{ƸU��%�"}��a6?b8[���3��99I:27���}�[J���X����1qO}��[�[+�XraeM�c�����[�R?��3��3HyC�'�t*��N�n�� (�^����Ў��Z|/���fro������%ZR9�����	,���pq(���&��x�{n�A�f�y�ד��8��htzFs�L�`�Y+��Tf(�'���� 0O�3�wʥ]�i�<t�e���)�3 ~!���&����ȨZ�zH{�8��W�4d���AY����&h��u����,n6:Z �[=]#ս\��
������ ����s�|#<O����i�w�==AV�t������݊����ߎ��@a6%�EQ���*�w�\S�S�� �zS�=ǩ��ʬ	A�9��r�l8�� X����I��s0��銉�J�t��8\���HS ��c[r����r��	l�^\��N�u� p���7W��u�g��!#ۓg-0��鑡4�J=�Ǳ`�qꐑv��Q�y<�թ\DE�^���x����s���B�kf� u��T� Y���t�$5h�W������O'��fN �S����$?��ǹ��q��ݥ�)/����g�L1�����m���|����'��$t�(�3�3P{g�'~���3W=�)��*�J����h��8�%���#z�c�q���_Y�ix��C6����@.�����B<4!��hc������K:t�AŇF	��`���w�V��5�[��Q=�Q��@@k\��%���6�3h�?PA�K��^��m�Z��s���؈���0�vV'[��4��O>�]�f�&�θ|b���WWyX��+ �����W.�w�����sP��&6�l�02�y�vue)����˓��svL�@w?|�pYf�t�_Wt���7Ba�)�tF���ZY\Ԟ��`�=��0�N�ǟ�,#�Ms��DuR��M��[�,\�5;y����T�Ty��r?�A���w2��g��^i# �cd1؁����!��P�?��jYU��q&���a��3��i�_�ў���O��C��JE�����;(�����y5J('��9�Z�Rsq٫81�ś)v�LD5|横�h���9/����3��^����N�'�gU��Q�6t��q�Vk92Y�onu�<����Ɖ�+8����p^�'���Ҋ�=	�u�lC�.2�$o�L�N���lRM��F[�vS��Ԁ k#��;0Q4��W񘾙Z�����>�S�q`d�g���m�rp�߫��>��3��'���>uO���9����c� ��p�L��'��ʼ�AER��{�C�=~��O��oV��$�X��.}I��MJ��Kу���G�<yX�G�?�_�#�-�����xȢ����z�{��>0�؉�\��:��gb~�╚"�* C �Y#�Q���˻}d^�c��=�W�}3Ҿ���ߧ��2���^&��#g58J���U��S{fB��I~ߣ�Ĩ���Nn��%�#j�&�ԡM�2>d��U�[ڼ�������jZAe^V�کk�Lr Y�^W��2o0���2&Ͽ�����4�t!A���5>������V�5�&7�!ރ��仮�oPJ�*1I#�E�g��!�͋,|b��f�~�y���?�%P�T�;�&>���j�;�������?���O}[����M�i��=/�3g���ix	�[�/I|�� ���Ddh��/�������5�]V���B4Y�2��C�����%��X76��������\-��:��3����}�u�~��m����U��9��5���o��	��`G��	](�u����� ���]x��B?]]�A֮�y/�v>sƵ۴[�1������AӁ�ը�=^�%��.oi�������1a6�S�&�7?��������j�r��( *�o����C��RK�W�"z:���J�`�4�}Ч R�vC�(qnfJk��@T�}Dz�=�щ���(��[t����m�>9�чG�aI�ׯ�9"9A"a'A(���w����\�g��Ê�ث���a�HXrx�sIͿ��ںz[ݳGt��c�O߯�ɓ�>�Ỏ*usM�M�0Xo��X�'�-�Gu���Δ���)eO�T�L�Z��҈��'�����^S�g����i`>D�V���Y�СM�)`J��6j�zI�ǾAʈ�j�������^r�9��&�V!�$��v�4��=�A�+˛a;~�oLZ��n�����<7T)���T��?P���� ~#GAY��Bjf�a���y��*Y��u
 ���N'[���jt����?���?��y�;���u���Ĝ�3>8����[���X1������h��i���[U䝜ߣ��}ꎏ+[U�����N5�я�;�Ws��S��)��Ef�*3wP��9�������S��>�=����Q����p�����#�N�UlnF��wi���P�O�w6l&=pZ3o��#Ӏ�S���Ϩ��K!hz��K���O�y�������hgx� �_ç�(~�H�{}�*���1�2�"��;��ħ>���(zd���ܯ4�03�n-�J+�-��0���G���Oyף�>A�CVZY�I<��u�.p�`��m�c�[����[�����,���7:���#��o~dv��sȕ �C�S���{�Y����{��߶;��B�(���}P�v��g�ah�Cn��7�zE�;d���
���5��j�)L�����9/b�˴ٓ�]n�oz�. A��тFJ���c�.]��ꆪ���\�m�l�61�������	��a�Q�n�D��Lt�y17�̻ޣ}���)u��Z�;�4$�R���C��K�ʰ��+4���Gߧ�O|Z[�b��Ѱ/����ʐ5�q���5Yc���A�C�2�X�A��
#a��k��:j���������D��@B#����Q���"^h&��+�S?�82|���o�v�y�O�[[�!ءt�K�"2�������F��=p���� ��ʶ6o-�����0���J_~^5�� #%dʾ���د���N�&;]�c�Ԥ��E����	� ��N��/���"uY��PQ��a�< �¬�h�$��F|���m�@>�m��ک�42=C��Q~�]�~�{�I���F�V
�~珨�����(_R>G�A�1r�*�S
���q�� ����z�EEg�|咚���n�+a|�� eo4�-W��|[RY3�����ooa((�6x=�t&��nS�fD��h
�p9	�[�l��ܥ�媖/<bdUf�>_��a9�*����-W+�pA��}/���]y�t��0��Z�0�I����GMF�r���#������=���ޝS��{51{@ׯ\�cr��
ȤU� �Vr�V����`�i��+�n�/��+�
rmú{O=�H��w�?�����a��ԍW_�@�dN����:Y  {�B`�a�szL����q4ah7i[.�Qf9R,��I�^~Y�\�!i����C�ѫϾ�&�-��'c.�[�?�=#����|XّI@'���_Wڀ��(c����+/����}�;�yۣ��3!]�
�T��Sj;���Ϫ�� B��yثw������jY�d������!��_zV��9Զ��C&�󰀁���X�����.�lĆ�ݡC����7�σ��l���]Y,B�\v�	C�FE�ȯ�uȞ'������Dmp�?���iA6B1?7���|x�u�L�����' 	,;�����]�G�O =���BO_�Y#s��aO��a���h����$z���-����m�qm:�ٟ��
oy�Ǐjh����� {r=&*��-��d6��~D�~s�d_X��z� �܏W��E�Z;���t�Mt+�5�ٟ��S��4(����?$TAzV��7Ȧ�6���v�g7���[)��x��W�\��Am�^&[�*�yR>�Tv]���9ʭ�-2/���3�z���z	myO���O����7kH�����T�5'M	FVu ����t*��g������6����⭫avi'��u�G?���۪���Q9Y���a�];�PR]�SY糩���;7u�����>�?�3�x�G5�������S�kld\+�E{vh��s�h��P����:�U1���2�Cڌ �:ͪ֯/i������<L��ӻ��яe1>)�ɏhqeG#�� L]7o\���-e�*y{Cم��ġ�����{7U����Y��Z�uK;��Y[����-kus[�FG�s������)��p����͸~f��9��4�5BmXL�憚���]���-��;�[�q��6�6���J?���4�ZV�_��	P�l��&,ޗ`�J(�|y�L�#Hb�Ψ\7�s�#��l< �XGw~6}L�?�"��^��6`�>��,,k�⋊Vv�9C��<���v����<"@6�9;B6����O�;t����w.�CB�����(74<<�A.y�uچ��_'F�:sVW^{]�7��;�i�|؀��k����z�Ň���Qz�Q���sa��c�M��K�O�Wm���SO�Z�	��N�坹G�;�{��`6�#���B�إ%�/^@�odܜמ�����N������l�Um��-E6���@Q#[����us_��Ӱ]�E�q���i^_Rq}Y-2�8�ǵ�� 8Y%���k��{"q�F| ���l�7!z��� 瀞��?�s~&��dg}��noW�tP�ݟ�J�w�h�x3��1��������M�.�;�ۂL@�4e�80��/�����Wav4,�x������� 2g��3�5�Kv	P��7�z2S�ɒ���Ub�Q-_\�{��s�e͐a�>�&I�1#���e~�OV�����d��ag���(������Z�YƟ��{��ϻ5���m��/����.�CYHƲj���'|Q
>�Ц���H����^W���w^W_�����]l�ݮ���͒��9��5*��X���_�mh����M���⮻�锶T�Ɵj`�G��TD� "���0��(��'a����ح�mi��l�(���?�������Y���
aQ��ԋS�J�4I���tT���ȱS��tU�[��qCt����ߣ�Si��2�<��W{{oj~����5��l�v�I�"�;MĻG��Y"Y����֊fG�����O~נ]�>��U��7�8��&	08`wkGu�A�-��*�~��`H�I�h%0x��  �N�p�hHC�M��c �X!����z����=�]�l���y�q �t���b~�@���i�+_�p��ڊ"��������5t�|Z#��\����A��6�Cà��3�j!�:�����lp?;����G2����3:�lہ 
[���Q�}�j�GT�a��@6VW���j�2@�������'O"�1��ͪSk�����7����cL�������ؒ��6x��<�L��}wh��X_Z��8�N��^�e�)m��R���0����T�Դr{A��M�\ݕL.�ܳ�loX�a`��526�a2 �Om���ݺ��;����Uwh�3�a��od���B�ݫ(�;9>�R����E�-,*MP�CJ�n*F��K,��y�0=��s��\�֍[�E��pI`�ܹ�d�+CB��4��ە%�/�E�Z�y�,nC3G��	;�>��ǁ�<v��~���!��P���W�9�L� ?i+���<_Hf���kyl�?s��8�u���p0�f����_��A�pn�_!��ū8qxϟO�����6��W���@�*�$� [h��=Ef�����Wt�O��E츩q�p{(&G�8D���߽J����R��RouU�tUO]yR�:p�0���|\�N�{�N�@˽S�����oQ�L^[�����`7��i�����W��#�%̾�QE��bNu��奛��u�=&_���[:��E���(��~(�V-�4�ն��kqKK|�@VS�H��­���M�C���y2�GA�%m����3 �"z�:��O�t8���gC�o|U��V���ۏR=�b��4�}��7�������K�ԯ(��Eu����G_Wa󶪰�\ǋ��(yX 6[M`�ٷ>��t�����D�=��j���kJ߼�\����U"X쾻������FƁr�-M��S��M���1B&F��MK=;_�FԜ�Ӂ3�t`��0<�y%������k�)����=q@��I�!�+��%�� �0��'�\_�)
�b�/�a�R�D^��~]�^U��㘃@i{Uiof���U�㯐yx���>��<��$ �)����u�41H�o�ͽ3�w�������u�u�	����Fa�CϾ����Sm}��a5^���|�N��A�������Sb�)��b)e �8�Q푵`��π�6��g����Q����羇��x9��҅�':{�%% ���R1`29�if�ɻ��\�&���Օ|&���t�Y�ݧ.?~����	��zK��Ƞ��;J`{n�W���ƕ:{N^�v��ʺ\/��774�gvM��ʫ� ��Z��8{J��*��;}�`H&D���>Ff&���;��K𯕍k�Mo"�&���1���D��~���ب|�b��%_yæy�K_m���1}�x�"�谶����D��=�������i����C���V��u��QШ���R���*]|I�nC�-���������.Ȳ�N���;b���o��]��A6���u�����=����0�6���3�#w�2\[	��붗��=�nK�i=�ol-��w-hf���L���֪�;ee�.dwJo�;���_�#��}��!�x9��H'S�$>�Įh��L�'	X�#���چ6���v�|Agy�L�yh3�]��Upd�������ČFǦ�mS��Um�Z��S�(=�S�����zM��B�~nD{'H��u-\��>�?�LTWվp^�|�HP�U � >�1���/I�(,.���@�J3<�b����~ρ�:�#o־c��?��_)��\؈���|:��O*1�\w? ������ �ӳ���;��Q�� v3a0�q'�@��Kʘ��T-nrF�X��6(�@)��ʏ~�(����k�V1�vRg "�y]�� g�`�5��VE�fK�BV+[���"��f�Ω��?&@���lM�-OAS�[a��r��*�(�7�0 [��o(� &<V� ��q����:�~	�F饭-�L�hdaM�?�O�=K�]��
�l�d0������c�.q�r��(��Ů.���	�m!��F^��CN�S�.���f���DG�$a�t)���(ϓ�>��aqK��pAɧ^P���z���qP,(	kiZJ�//7M O���h���;8w���P�5�8�7�Y��l�̞o�L��Ќ��3-�b���J�!=w�R�L���fҴ���
��Swx&z��1�����~���]H-��s����}�T����,A6_,�Um(
;�U,Ԑ�s/ qЄ�̐A��W�̏������^7v�j(:��)���]�۫r�A��#�f��WG�w��=�Y^}\��ɺ�sG��<���"����Z2_!���#���Q���%a)��wK�}h����h�{F����f=�ޜg�N� �#��yb��_�{4�N����}���bw��g�����hV#� ���������N=���blI|�c���;��zh1e/�u��󃯛���ݧAg��ݧ�����6,Y�o�$�%��D7l�J]�����+���f��~�3�G�I����{Zl�a׽oqY��?�QK����W6�5�X򙸲|6xl�Fv]ka������~/��c�DabR��F�W5x�;؉W���nD�|B��#�ܧѹ1�Ȝ��2؅���|L�[�dS^iG��Mw v���+�l��#L0#u{u�G2���/+q��F����K*�OT�ܿP�?4���\�\��#�;��X���O(11f#���Z����Ͱ�$0Pw�y��'���ft!�FFca����#E�7�N�F04Rg?z�Y_V	��T�չ�wT���b0����W��8��k�����Go-h��5�t�RW����O�&:Ȋ���StaI	����H�l����`nC�U<=����^gJߺ b�M�A]S�\V��_�j��׫�vK=��!V����捱�p�����a۱pd3&�爜�:Ƈ����^)u��q�����Bvc�s%�$�H�U��2�9(�a����|�b����*/zg�_�����흋��@h<����S�&�lz��D�0���~�^ޅ�=�G�ç�ݫ�m�����<l��Vԫ�^����F ���럏O��*[d�u�< p���x���_�ɴ���t`u4ŮV.=�O���xN�vy���sH��(rp�L����X!p��ʥqL��ܐ�/�� �Ml���2��9����u�{*�&Q�{���g�l7hv@6��{�K��� ��]�{�N�3��iE74x�E�~AS�K���J�U�_T#0�"�]��A��[?�_V�<�l;����%�EDgy���W�/��_��Z�����`���A�D���m�=t��ƶo9zM�u�a�F��C6ҍ������{�#��"���~�`�R�i�s���r��;I�O�i��`�v�7<l_�p����4p��[�@1�|�d��j��#��D�h=�f��>�U.퍊��I(���'$�?;�Z^Dნ�&Y��f����o�T�9\����^�.j�s����6>h|�5 �|�7�ѝAY���0����G��ds���d����s�^�UG�(/�����3��®/',QRriI��_R��;7C9��w�-��xH�2w�����2?�)2��J+�������W�~����!�X�����h
G'����/l��08�oW�h��$^�kz�f7E�3Ś���(����H�4D�&�l�.X�@!ago#��L�@���p����˻��~@���׺)����f��yOHzXV߂�!8x�~����7y��|h�kC߽V�'y�_�L����#��Մ�JxϾaò�����P��7j6:��B�����"�8Fڹ�z�)p�#)�]c�Tۇjۉ;8#o`��t�W���`pL��5�6hOX�ְJ�Ϛ}ڑ����n���&6��'��.A���a>]�p�6�wpi�Swt���4���M�Ȫ�"��Y�^7'5�T;[�z�D�![��Ďh��럇ᇶ�ԝR��A%�o�|c20��aO��J%E�zp��#�}S�ާ��M�H?l�	��5Ɍ�/����V��������U����5�#�>D��?��s��㏫�ʑ�@�ѻ�4d1�5�l����zlxr;�j��$�M�����%��d'���M�kxt�0���/�!�T3K�Mێ��y�	�zv?�U����[#P6�*%�^�ﴻJ�ї2l��lP)Y f?��a��Y0�`/�Kx(`�d�I�m��~?�F�=�m*N;L\l1փ�м@�[��mw1�I���`g&����cn/ٓ�7�ɆN�t��ʹ�/�ٞ��1���y��]�π%|���0<L�����y�:w���2��g��1�V�Y�a��~~��j��z��r���k��j��=}N��>�2���k�RťU5���h�r�>�uN�sj��QM9����n��_Sّ\�;8���K¹����z�n��.���_�G)�%�d?2v ��=�����&R�;�]����'5�￢��S����������Q�UXL��'�:���: +��U�8�j�Z����D"��D:�`0��R9ս��v��VL
�(Ej�`P���o�㒪� ����a,):oyrǻ\� R��S!O�x��k�`�a����roth񙔭�ՎE��0(ֶ;��
�����h�5�N�p
��1�70�����D����f@��"��s}���$�YD����v�d�|��{�a��X� @��<��4F���o3����X}gMfS��i4Î[/	4�G �m�:.��]R�n���"'�f��&`((����M�gvf�:�tgB��N4釙��أ�瀗B��F-��� h�A�_	�v4O�wzd��]��������A0\>��J��òu�{ �W�_~��$`�b\fݩ&�C�t�3T.I߰Q��u3��R_l��}�ݝ�^��⸈`�;8�KoxIj�u)����r�_�iй���w��:��=�󑈱��`����Q|.=��f	�%��A¡4V-�{���c��;�	�$�c�@��s�4�	�Av迃���������d �0<h�6ז���\��v�m��1t�-��"ؾ�5-j2C��rIg��/�#��t�WGoY�l[��ՠ��|6��K�]�;M6H����:�p�g��j׼d�>"�4�ѻ���UJ��iaWس2d �>ha��z����{�=��� ���H�����;
���P(ʗ��ccؖ�;�!0��jaN�"�w��|��Cr{��h�vЇm��d�/��
w&n�?%h�}3y�Wx+������.��Af@�m/����:��v�v7��|N)�����_�vI�'�A��@U��IoA :����X�Aπ�R�DF���hU[��t�HC��P�3V(��cݮ��P #�	4��N��ۀ�GԪ��\I�����s�z�Z��̑�6�<7ЬxGg=��#�yk4���� b����ώpmLw��s4���p$��k>ػH��`q�J����:�8�A�<v
8�NJT��/��aPi�f!^edFn��a�l�T3�|Cn�5”�WN��+�W�xvllH�I?�Պ��|`?�����tQ��+�U�D3[���LŬ�T�j�n�a]�}w�����\ء��g���\!Pٽ����3����q�N���h>6����Ȯ��y�U�;�}N��j�O._T}�{y������A��8M۽�^���S�d�G�{DJ���a����5��bCy�2a ]J4��X8��և��\���*�&7��@�k��(�۵�S8k����w��ø)���Q���>Y/��N��䠞�=gc��E�3|�{ؕ<�Q(�P����+�[.�0h��8�6ީ�� g6�Ju����|�0�f�-8�~�O*��*�-K�
yW2��~v����_Ҡg �] 8�����i0�����aG��w�N{ٌri�W��a�^�#KLz� ��)��~��d��g46�l�Z��~���p�Y(��w=�S�b�J���|�6�B5�(�NR���#�E�!��%������ c�`����#c�g�ZC}��������`��i{k�|0��@=<>���U|f ��e'�z5ߖS�Id�V����r��
r���2n�}�d�C��\F%|2Efjeb�j]�)�ҖA���}�O%�	���8Y�W!��$5wv�����-���&)�^%�$��:���/*3�Š�� ~cuA�����8�Ǎ�Q�R'�9��԰��z�Y�Sc5��Vָ������&������ * �
�m������Ζ��#:7PguK�Ʀ��n���ƇI�FQr!|ֆv�zNԮ�8]*?"t�{���;�Jm �È�|��jUE12/Y�{Y  ޼u��ˌ��i��,����c����_X��!��|� ���(ͧ59����\��}�l�:S9;k�"�`�F�qڀ�p}���Ɓ��3aج�lT�{�yL�hl��|;l4J �7`�Q;!,�N��I���>�h:��N;O��msydRC2^�Qs{���q�����^���1�V����ʎ��>��7��D8�k�C��i��:�%�5h�� ʻ{{��oF��Q�ob��Zu�͎a�f~�U��3 Spz�Z��6�-oo(�|��PB]� .�����e�A�[��졐�1�q_o��oR���M����{ W�`5Kc=��>�!�<7�����Ŷ7�yA�Ss@���?�Uf��ܰ3�+Î	�I��`���G��.I l�O�ň�B�
�)��5�a���K g.���XU� B�L_}Y�	|�����\��@�9� �7�h��'��W�.`c`��z���]�}�lq m�����@���q�,�l��;���|���a��ǵ�\t�O�1K��w���;(�g�g[�#�n8��w�^�9�_�i�'�}�KЃ	��CU��>�d�]��
�s�z�Ù�o�(�v�V"9�**�Ż��}��� ���f��M��r-)��R�I�������\�}Jy%��̐��XdFG(iuV��6��ͺj�G X���7��è�Ð�q?gWj&JIhێ�5�φ�݇���)��B��    IEND�B`�PK   O�WW�.�ɭ � /   images/946c31b1-53e3-4800-acb1-710e2b91d3be.pngl�Sp%LԮ�ޱ��'�ضm�v&v2�Ķ�c��3�m�����N���U��~�E_��^��%I$x<x  �$-%�  ��;w�B����������f���?��� ��ލ��c8')m  ��7pӂ�󿤱���������������1������������)���')���G��������\�7���X�/4~ |qI�	�y�x�[j�o���o�hf�5_�r��!B�A�*���͐b5RtX�@q����%1�A;;��&	HM!T!ؾ�ǹM�4���'�޼+?Fֵ�{�W��9���]�؏|�ڏ65��[��֢v��F��7���W�b��ΘXX'�A�'��ɩ)Ó�������ǹ肭��վ��uu�^�C���'��^^�)�!#5�A�s��"/�o�[.�&�8�B��vg�k����)���_"����4G=�-��JqJ�em��_��D�[[ZM,=8ehG�EM�j��y���1��,9���9k��1,�j�>�&..kJ�>)�-X����Մ�RWJ/j�F>>�KOঢA���e�a�Uc�[g/u�橚��c��P0���)�`�g
�X�����c��̋Ε�[Q�?���$S�\������Ҕ�k����nk�Mѯ$�%��0��{:�wկ��n�z�|_*���o��B���zz���TQ�I�EbWK~݅=k+*�)e���H��0����[�T���"�J��W�{-me��,��[���?��v������ؙ��g��#����w||�^���&Kq��be��Ⱥ�����5=ΓD����"f���T���A��SE�Y�|�%H\a�ǥ�B��nB��(�.��Q���{�c.�G�����>�~����e���xxi��7���ߟ�_���w뢻�y�2��f��v����9�6�D#Z<%�F��
GR�D��:���cFE�"5��^_;��:�k�c�o����Kke����v��Sz�6~�������C~���۵�6����=�MY��j�9��;zO�\�ޯO�֙xH>�ta2`Q�Z%��cj.��5���S��zWVG�9�ԦeL=0.|�]@��hkË	���H�⿻�Bv��Ъ�N���UUTDڳ##!T��=�ؐ1�O�	�2��F�V��t��+D�P|r���O�m�7��;F#��$܈~A���p����O�A�BX��N���f̾@c,���`��Z�S�fTʠ���:Ma�n	�r�V�G����aУ	��h-L����M��>�m!�A=#��c��3,-jT�T�LθZ��/�£�<�s:��LJ���T�y��¶9����g�E��dgJ"�U@�+GS�W
J�n�R������p�?��9�By��S��O�'J	:�ݧ�><���<�@8���&2Z��W��P��w��=\�ߌ~���ʼBJ�uPK�HK����G>#�&o2��¾�*�^Vl�^2C(�=g�*���+Ī��W����v<���1su�4��&u��W˾#�$��U�g{ܦ��`W)�o����l�3�G�G>E�I�
�{DxȦ�GV{�Z~r�o�kz���:z_j�{���i)�k�S��<��Ӎ��*�9.Q�ˢd����sH�W��	ĥ��D�?����y�/��eD��}B�̀�dᨇo04��J��|�:3���_�YY<i�x�������r�k���=Oh�9MX�j��b��VQy�|I�<,f��CJQ&�P:�j�s���SH?�|T��ݚQ�K@�?�VrV��L�ڏ�Hd{ɍ��3��j$�.!#����x1=]}֢�CB�0�W�2Mx\��l�xFz�%��/χ0��z�C՟܈0V_<�n�v�2[��G���x�C���+�ڝz��_''on`̥J��۫����f��7��R��LJ*Œa�ti�eE˫��4D�g�]e"xz�Hz������9�+i�����C'f@��2�/��R}o/ΏD5V�~ϲ��7�h���.�C���������!7yPP:N�6��GD(�}�����&�Ey��_s�8�j��tt�/]���tF��cB<\��Cw�!���!�RZ"W�����J��G���x���},�QB��B�v���1;87b���=5շo�ޏ�l1s���đ��͚a�v��7�kn��9d����o�E���P?������x���C�[��N�������M>������$��@��iw��~�/�ծE��ֲ�y=�9	w��������W�
�.����6�/��&m�+
�ُ� "�#jhjvn��f�6-�{!B�/�Kv�m�$�K�bx�.�OǗ���̑��jw��~���FJ뀑B�<I+^Lu*�z����FB�խr��i���c(?)�'���P�Ce���n���j���5�lB�Ǿ�"
�ҷ�@�t�C��|�w�@c�����p��!�T"�x�����x��C%���NG������A�T�2��i��-�N�t��G�Ý�6:���he0��&��e�)Y��K�����΢��4o�?E��Su&�����ă��R^��:���g6V�r	�k�0��'ͭ�3��$;�:�/��c��zg��Z�~�-��L�[�����ĨHBd�koSS4�=��q�;V􈿭�(�c/��*��-�c���7��_��?�@I���;B�,"�A2W�]�6�U�Iބ%<��4� �!�l>�4�x� )I����Ui2��/ic��I�V����C�[����[�����v����-Y��@n�ߩ��w�N� 3�\���7e�i#%r�5*� �	ơ�Y;��U)��0\,�(������yYWA�?�SW}ƺ�D%L9��>x��Z�2+,P[����|40���^��=����8����bUt!ޢ���F����O��/hST��@�	%'��	�m�4w�E!�3�f�\�<y�n�<��O�bљ�� +�߻^�s����R#��b�!�����Ʃ=>��#���U�urdU��e�|+l���z}����/q�яӚ�(P�����\�P�%�IQJ��������^�ӊ�<%��T��>��8��xJ[o���b�v�K�aP��OL�������5�_	���_W^v��Ғ�q�F"0H�v�)�s���[R3n�xND�.�M�8-����݄!���[�4�]2a�GtKSC]�xx�O��'�O.�	��ӈ����P*?��N�z� q��6�;����,�&Y�������oN'3��N�_�9�����t�e��4Y�Դˡс�LV�,���V��P�
G��5b:�|4�������l��H`�V5����
�AK��/*���cb���7��>�@��qD\���(*����~�����GR���@�пP��uS��-v�p,lVȆ�ʇT�T�F��z��3\pdbx�������ٗB�U�O���/]�R/�[S���]�?%�Ϫ�T�K|g�mX��qI���<%	1X�I��(�� ��xdZ����Jg�f��m`V��i��ش�S��gLZ�z/��~|z2�a����Pcbu��H��������|�72���c��Պ�Ԧ�8�{�<#�DF`.���PaW>��B�C��ԡ���J��b;��������=�x6�%�{3y��NT ,�#�H�
�#r>��u��h�t�KLN�
O.'�zEk�,�_�/}W���^�wB�31U?ӳ��h%�u�o1��{��מ`D�rJ0WYpF�T0VYD�5k�?�wG�'���Đ2������i*uK�f���H��8?4���o���h�Bf>��c�a�䁽�N�]��z8L⨞�uI6��R~`��!˻̉7UUsnu�%,�V*�m@���j�F�ċ��O1���飫�����@ϐË՜2��j�J�S`��m��w�q��'��-����ab����^���j�PGGeH��}e}�"2O�d��YrPq�7��{������
�	e�^��b/'��ێ���ŧ��J���z���%�d=9�,��p�JtY�����|�%�7���缘�w�O�����$�_]����� ʦ��f��1t�mF,�>�HE�7o..�%d&jx`�ft8E�H�HG(<�C����J��cpo�a��6\ح�1�q��4�lb���y����������	�CeBPOu�8�"Tb~Bw:p�#t�Ȭ r�@�D�>I�rb�u=��|�,�	[J@��55�����ҕ�E���o�~��;���\�Al�:�K�B�O�F��踅A��lt�a�������P֕���X��(0d���5z��~z�\��ܬe��i𡌈�8Rރ�.e�0Z���1TUգ/��3t����h�.}�n��i��T�	��	�H�)��^6��[�0��\]^�\���3W.؟�<��<Ґ@����҂&$_�//Y�&��,-�UP�Br��Ñ�j$�����d��M���"�?xv�y���U����V\pm�K~�����O<'���vX�����A��Ŗ*��[��8���m	�P0k���n��:�:>)�_Em��)bA�ˣH��@�����U�c*��`+���"���M���}d΄��D��,5��ywͩI�a}j��+�������S�0��0+K��1۱�<�gm��e���7y��q�8H4U��0�b`�+��4�/����ڼs-m���8�G�n���bE0���nM������aJ�i�@���j�+l	.�7B�c'A�6ZR�~��z4C�p/j�cZ��'��z�--��� H�'L&(3�e~��A��F�~��N'���gw��nfmc"qr���U�E^�����jTG��{��g�����r���鉬X��8�֔�������9�OMI�2KJ u\��\m����F�1&nb�rcK��[Z9dH����8�o*���QG#ik����^Y�߽��$�O��]H(H�X�{W�iyr�z�t�z� '$����v<��9�گك���~��.rG_�J媟�0��L^�({�=~�%H]�N��Ί�1H�idd��#叮>Pӊ6bb�^��i�ľ6��|���f?g�T�d�x�[8ѯ�q�Z��4��&��1e�od�|��z�W���Vl��RQ_"�\n�w���/��.NԀ�����#�𝙛��/�Ϭ�-AL�~���}�q�嵕q%%�e>�Ic~��г�3>�����S�CA�փ�`4�IU��b]�XΧ�ת���VU	��zP@���e�ю;f_:��Hf������ߓƮ��+
���R��n�H����p�N���G\W�GW.�jv����%/#$�hͤ�����!YsЗ�qԐA��_�U35����O �5=%"�Ҕ)}���t��9<l�xT������/.��܀G�99���E9�ء��gR󚢲����i���Zw�Q#N�)��9���Q�9�h�ʞ*g���������t��5P{�����+E���w���]X��b�/�r�v�}�Ki����Ύ��[��������� �䵱�� �[[	$'�j%iᴙ�/-H�j�sl4R Yn���1jp\k����˺(�K5v�z�$|}Ӡ~Bau ̩G�\@K@���b�DQ3�Qک>g�VDۂ>���g��$�ʜ[!�k��ց�z�>�l?Ġ�ʺ2���N	���߼P��+�d�����"d5�D�|��7��-�n_�L-�_�� �ų�j���dt���6ڹ���;ힷ7�4���
q>}��#Ł�6����;S�����'� �IU:�a�!$��l~� 
;gC\M������ncg*�B��2���-���O�F����!s$����XXn(�F(B�J���+���Q�}����>??��ƣ8�<�ws���l֘���Vg<hn�97���C�+����r�������8~�ϴc��2y��Y�/���ͅ������h˼(���8&n�������_��DWQ��\O{�0_��#���a��{���O(�b�G�h2�S�9��䢷Pc�p���Z[LҀ5���`��hȬ
��H���!�B7�5ɘ;é�^�EwxS�J�xS��,�"w�␲��}XJ�V ��˹AV�߷?lI�D<�MA}�N��~�fF��|�~?��']b߶�i�OMO�b�� j�����bc�_�&[�"5$����4���(�q�X�����N@E�q�.�J��w�M�	���A<Ɠ���0�Xہ�T-�ր����
s<��E�R�s)�D���?8=77����A?�V��P�Ϗ���`+@|�}�}|�E̋��<��Gu��D#�P���)M��Wۧ a���u�{Kq�!|��x�p��&��k��斜T�q?�Ge�C���BcO^5�����+�Sfnn������16��_-t���͟��m2��֤e� 
��*�A�M�(mqo2X�����6+���-H0�w�>=�d�#V#D,a���8Ξ�bV1=dPI�{�&��l<��i����K�qm'�����q�Y˄ cyM���Ė�Xv�����jH�4�S�Y/A���	��l�7��!�^y�%�d,���(3��&��c;��$Si�M�)HW	����)�%"j������:�J�R��(쨠���5b?��}��BA�.�5U�D�����{����o*�|�@��_f��^Oz����#C-M(��e�$/��E�"���'\�EՀ^���=��#��id��<8�x8��Ns�c�@C����)�jd��� �*ВEcm/�� dlq��|y�=7��'�����#q�\,�MEi$��(�xU��8N��O�[0����1�EafVF��yd��\='��O;��?D�ں]J���H�n\�$R���񵡌V+fu K��W٠��\8�O��^ˇq]�F�Op�<���,���{8�.㞡�����m�dZ�J�`ųȯ�F#�~��Aa�G��v��m�P��	; �g�Kq,ܥ��BZ&�-P�2R��
�|���{E�IW�ap2C�� �!��+(G�&�c �����#�7�43��.��2�U�t���V�6��Q(��E��jb����)��8g��V6eQ��3��t�[1'�pտ��4��?9�1xAo_�zW�ǽֈOQi0D�}k�L��dƪ4⍛��_�.~��������vW����JWObqZ.�(}�F�mgc>���QUF"Yܘ`襭H!����
NJ���ѵ�P�e��C1+w��:���ۿ��t�Q�ۀ*AP X�E(��b�FB��m��$�f�FZ�"�ʸ�y��#Y���Tp���Xx�"�!�[���ɜV#�(mSj�J�Od��L{d��-���µ����d4��P�k��&c�|\|_h��M���vM��"N�
�~jPJt�T���dV}��Q�\b�Gw����Qȍ����<�1�i��y��v�ֱ�Cmt�j�@���{:=˟ᙥ�\�
:-�xQ���i����
V�u�=Ou[����nXs�t����&<u��=�⎠�c�G쉤0�u�fY)����|sȜ�Sm���H�F^��R�"W]��'E�G�M ��D�"�"�
zz����t��i	N'�S 	���a��2g��v�z�������5
��nE͜x��Ӎo�\#�9J�FY*]�_l�����]M�Z;�����Q[� ^��1��6-�C/�!+>��������y��ŉ{G�:�.�x)����#;��o�����))�����U3���g_^Ĳ�PӜ�^�f�<0� �A�
aEa�F��Ʉ�:+´V��3���6�NR�C'�Z[�l(�R�*���~�P陷e�q���3W�yD�1T���i������=�	&#���~/F�D���)�����3�<�a��/i�H�БÑ�*���u���O�]�<l��M�dI���Mb���=;�V��t� [���:l�37����B�8��m��u	�|�����t5�"���˘y��n���H���>#e���H� ��:{{JUY��>��<��B<t�L]Q�~��U��,ƓŽ��uDR���L����G��k}��,�X�?�5c|$Cn��j���m��:���x�/��r�~4��7��}����HʴZȦx1/���&$$t�ݧ��'$=������KJ8xxy� �u��K��͋�`�4R5�8{�JHX�����]G��%𙭁�Ǖ�+S���/Wq���s{q��ij*�� KR̟4#�*f�����0����[+b;3�8�y�g�����K��bю�2��4�&Zo���)$Fh�(1�i�l�m]6 ̬��ߵ�*ύL��k�Z6�D�V�U	�:xu�F�\�n��d��M�N��OcOWy���8>�~WܩI�tV���H?�O[EHN�b�����X$t��Ip�g��@C!����^<�D��y�������7�|H��-#,󁽊S7��e��I>sZ�AR�M��zE4F�r�Z{�q������nwW��˽�fۛ�F�?��9�3��:B~O��m~O5'����k��b�-t����z6�
>/~�L����|���@�!�Z����8��v"KaW�����f䴎k��lg�,k�ͧ�c������Q���$?��\�}eG?4<k6��u����P�cwhdJ�����*zh`^ȮfR��&�M][���]�Lf�"rTP�q�rc�]j�^+��A9$�c�l�S�ה̻<vH�\�L˧�����]
�����������J%�pE܎�XL�`���"G$+r�2.��G��N���EKE�g�p�����K�_#~o��?�K�|:}��ޖ[��� .STg���V�ΫB�d�&'3"ֵUfD�V���K�Bs�X�u�&3o����uu�&B�d�N��\��y>�eff!������d����yt��x�e`��<�|l����1����P���z���ն0w>��8��Uܹ�·`.�V��e�6e�M�7��k{Z��y�R
�lTv���&��O�C�0i<�h����&���(E���Y�C��/vXm�n+סr���=�n� �z�q�v���m��&��c���܌܈�4�0���r�?P���p�ԎU�[c��8�iDh��3�\��K��W�xH����p!����l*��)<4� �+ 6X�(�F���hlll�ϩ�D!�@�ڪxr�ƀ��qǾ��X��r�
W��Z�	-E���:��d������F�?�)\��Q�!:s�!\`�&�%a�'�ᛗ��6�	C��1�gg��y �����c	����̴^^��oA����2Yu�̋6kb���Y������&��|W��ϔȎ2�l�{�Y~�c��{m���L�X5f�dw�Ɂm%�sC���_��EQ�-ۤ!oCt�VF���B{/������mĔV#Yv�LCW\h��X�lװ݉��c�D���r�[�˃r53�|���h���XrQ�C3�
77/|��r=7�gS�c{L��f��qhvַ��Y�3���VU��Bn�^ZyeC/����0�@��{��ߣUm�	���;�z��6����+{���-�J�C�`0?\"D���)��:�.h�Z?��rܦl/-��W����zj3C]m��r�#����F����=��;�E�}�����ڌ��E�O}�F0�b�CZ&����ʎP8�H��?H=�͆�
����u�;A�Ls����ב�H��5���<����ƍ���}?��*�?�s�KczA�)|�deg���+�_�ӈ&�k#�h��=�uW���>ęx�S�<�r<�����6�7/<��>,�15M��3���Za=KD���*á����aS����P�־�����l��hg��+o<;~j�*B8<�dhS��1��ێ��h���V�ȷZI���̇�\���$��?�N0�����TW�C�AkL��K.X%}Ɛ	�ONJ�FK�墋^ɬ}�����"�Q���բ���⮐�2��켈x����Ʀ!)��S�c2[�o�3��X뚚�0�FQ�1�ί_/�zd4��aۛ�[HVL����XQ����LѦ����qM����{6�������Ө)��=�\�dɳҼQ���ʕ�Q����GA���c���eݱ�ϱ&߇^���y�`j�!�h�[]�F��� �*Wd0IR��/��e���dR��[-ǫo/'�̴�i��fƀ��0�e�A��=�~(%<������ҙ@_����x�QC_ų��c~�;�*�6w N͏%L��z����U�������Օl���r���	�~��R<�+�:��[|X؁�Z���x�R��.S\���m".%�ʾ�J&xu��F�EW��I��O��\�^'7J؟�����y$���Q�M͞.�"լ�N�T߸�3Eܞ�!F=��g2����-�၉���)<��	X@��{AY��Z�o~���D	��i�2��s��|�ؑ\+4HG6G�b�c��+l�QB��F̈����1�ѵfO��,��E��#O84�+}�a������ƴw��P��0�G�,��3�suu-��cj=4'�\YDwt^�ꁻ�<�]Znu�[��O�����2]
�U�|�̨�@� �E���9��~eS̺[�-�~��< ���V�3���siVr���;�si-M\��ft a��CQN���2m!�Y��X��oR\�{�e�,�k�۸��@�o��<Щ�[�l�։�Ź��B%3���zR]9����5ϡ$�ٔ���r $�_ڌ�m<R�`NT�'�>��&�,��<�+�J:k��9m���"^���?� �2���W�k9���j�
�V��e(����ס ZF��հ<��J�L�a��s�⢟4곡�I����%�yD|��Sg?�������T�}l��ĕ�{��9�f��٥WU��'Gpc&���d��ޤ�r�`5�_ĭ�b��h_��&��&�-�$�^���Z�9-� q��IIf�P2n��YYۋ��������d�]�4�z��ඒ�̷�8��5*�괷��)�'�Z�_���0�J�M�w�Gs뢤�x���v�z�BYu�v�[5���.Zg���;��h槻>f<�H�m�V�)�ݍvF)��<��D��y��F��+$���G��l�H�1��~	E������Ϻ|��l>�nd��oiT�~��#��u�i m ����+�"��t��g2H��Ƒ�2Y�$U���} 3y�����a��k.7"aM�W��Q�a�Kz?B1<�wG����vv�j#��o����z�-���@z��W>��B�Uѽ�+܏0*���8���#ׂڮ�����sqX�h2%:Bnʃ�|('d>��џo��B�����W��)��al�g���
�ƈ���ii���|�:�$Y����c����J�����
�{�s��T�4��fh�=�A[�V<����9�`+����X �mu��(����nX�kX�ĝQ�?3K=a�a?k���Yi������,�t�y>����+:I����Ŀ�-�#V�쨣)	ќp���v��OcdJ��93wI?���q�J�a�ބ��A(����m	(�S�}S,1�m1�RU(�(���!Q�g�Q� ��7%��"݆71�2o�ה�I�^�G�^��-�x
�0onx�&V�f&�e �w}5��?��1
��e1I��ʉ��'#;��Vxm��"�^��������7ע˝�=�E�yE8B�Y�����8j��mŭ��㶊�&�Ն��h}g�w{>�T5�d17/e��dɂ�ׅ��LbC)[��F;�p�e�TU��\��J���y���k��Rj���9"OMa��[?�ZT};��,�|]GkК�|UP���cX��'b�P�@�����)�
MxX�@�pМR<>�8Sm����M	�q���ȣ��,�9���a�D黮�R�Wu1b�R�,_wuK�b]p��~	�>3�x�!!q���_u>]�^ua�?�T���4�����(���qą���+/���3���Kd>$HJ����8�s�}�����o�<�V��*�/���TM!��⩩�祹/�������{.<��=�����$>N���������q�/oI�,D֨M(��l��/��k'�3`��������8�,�3ͬ�w�����3�-��R��(���LY�H��<����lZ���Z)E�-�v�)A���;�lW����@ �<��ler���g9���P8>�,p	�8�ϖDc�F 0����p17S��X~c��py�"�s+��+���� ����H�'�Jb.�y�P;CHr��W���%Kۜ"rt�+c����H��Е�7Ul���#��d*�	�����a�z�WW�5��kgkG������o��Z����v��t�tM5C��jb �����6�
�C�]˦�uq1p^�	���/�����s3TB�w���]�6����� �љ�u�[F�^B�3������ɜ��m���%�j�:��#8���Ѿ��s=���JX.Z��q�~,TSEd��uN���ʂr��ђ;�}^#e5P�lK+'iX�� ]�[+��ϭZv�+�B� :�8�E��A�I�_j?�V��b��ϙF��N\L�\�m�?�������4P!`�q���b�PU��FA��$%#��
�-��ڭ�����96UHd�Rv8 r�g<�{Sn�+0��n��K�v�R���z�V�a�>a�p��Ik�B��j�W�L%�a�"~�Ū*玌��*��}�\�/W--lme�Y[���#7:7��������Q^�"�)���)�Ӛ 6^o�j�~��R���}�硵��;��0+l�)�0��Y+�):����6;��-�搁{s	w��/�G��[)�f��Lt���9�)lMhx,�b�D�٣���ȯ+)! �`�6D��h���.���E���2|�De����Hf�D����Db��Щ��u!��YRlʹI`�͑�u!��9	5��
�\u���	�_�����n���2��#�\/�#�����("�b���@���U�JR#�oե�x��@A4A��s���u@�J�ʨ�Ũ���=�\2�����!��I���;�N�W��I�5��Ā�UP�5-�ϳ�v��T��렺�|�����%��8������6�<�U�W*�s̸XHOmu,Q2Ѭ�ے�����F�Q�jR��xP�j�r�*�F�pT���8ݪ�c�OSg�����RgFIz�x8_���D�^����X�������F��Em�b��N��E�c�옭�k)2ڪ�[8 ׃�-���{�&��)��ؚ\.�[������~z8��Y�y�Hb�A����VM�=#[v���*�Ŋ�%lȺ���骂1?8�@������ H��Ba�@� �2�l�_mz�U~5�0������(�oiqt�r�Bow�CA�V���4���n�5#�%�.��fJE�3�93�,����+��P�v�C���/Q��0�<���ܩ���̴��h!�4Y)gU�ɍf3��O��Y#��ٱ$�(��q�o�9�=$*��=�@���r�������H�g]O]ʣ�v.E�"<c�GbſNcq���o�|�̞J]zVc�,�Iq4w#�����Hd�j��²�a���Q�uq�CS�ab�M�Y#��i�Ө$tG����>�D���G���e��)��}�H��Drn�:P{�����W<A&x��T�2zsD���>���3�s�B�:���s�x��V��0W�g��h��V*�Q���븈J����)�x�~��o����V�?I0��h����u�3�Q��iBrUV>wy	�N�N���������O������x�&4HJ��w�ջ�UM��բ�gM�/�]��}��7#�=�o���	����G��[g�����,��g-�+�r����̆�5⡲�1ɯ`.r���o"��_\P�%T�&�5��Ӕg��e��5����K��H|	!�[/�0fG������΄7k�F{��q���by�����V"2���b~u���G�L
��~�l7�ͩ�y���e6ПV⃟�[�?;�;�2�;�/�i��ɂ���+~��z�` `�Q|��:K�=�5'�5X����_<-5���دg���p���+:�z�cZ����`�/���R�=Ӫ��:�o}T;B5�SY2M��Y�� �����X�����a��cϋ_r�0��/3DFM�c�c�O�s�"�.K�̏dH8��?�vF��9�*;P�OJ���i�-t�Z�^^����?r��/�e���z2���g8���(��1������Dbo�pN���X���5����-���eH��k\�$GD�*-��0�R�V�F �%c*=�Y@ ��)����Ez�>:U��-MJ��:�6�Ł��,/i��@� �O���(�vG?~v���|v86Wr9�1e��x���?�����Җd�N��i�7�N��x������2%�������P����T�}f�6_�5Q�u�YV�0��K���3���9x�0Xe�i�j��G0e+( `�d1,��|���".8�����1�-�H��
�b%,g%�Z!����%ܖ!�]��Fr��p��S�y����z ��\��p`*k��������xz�jF3n�>d���ߞ��%&
j�M�OCSij�S�W��.3��F��j V�"��m�=�����6?-��R�-0�����Q�G��*�Bà�=C���(d�$�[m�CT�3��S���ԯn�r/�J���J�?�FC0s�Q���>�O�6P��|7�@\���@u/T)���x2u���^��vK�:B�A �:��Qݰ�G�O+~�4�>�������q�{j��P�ڣxg��Go#Xh��A[:�$l!��#��ۑ��@��P����,���R[�X�����d'��8�I;���.������R�'��xtt�����:[��l��f��rU��'��iG���)�;��ݏ��"��QT�T�6yY8���8�f���(�Jf.6<b_W�W�܈\���37mONL��S���\��΄�>�R��ɘÜ�^,<:x�jj_���#�/ۘ��*,�Zt_V>tdS��^q	��5KǷ�W���e�5n���ssފJK̡e����`��3�d���ta�5@P�����ϖ�	����6�Z`��Z�h�/d��������^睤XT��>ja�w��`�Jv�	T!���RY���J����I�_��!g���!4��)~W��ۦ�8=}�#w2/�d�Jg�o|���0*�VF�&ZY��6U1���� ��Uc3�~(N�s�����ߑ��;�����N��h�*��<Ddd�~\%ґ���'t	���{A�������1���.%��A�g�"���O�#/�M�W��y��%��BPy�?��/��#�R<Wnyf'�|��B�a�����em����S�{ 7�s���!ɧ� N���Vǵ���u�;��`Q��J#zR�u�9\��!���	�jm�&�����=�)�a�m>��CoA�2\1�u
������>�@��g����l�mI��
b��z`�iDӒ�̥��&������w߆�:��U#����rՄA.C(��0~��U3�{%��m�(��zM4V�N��:�(|������n�%�ku��j@A
�&�{���p�v(f
��ר���v��`�{���#y��#�Ǜ(����G��y�1<��3�_�q��N<j�Ǆ)F��N����n}O�s����v`D۝�x`�Kw�Ӣ��|��F�v'-%�ǎcP����&F��0���O�P�"�|��~GUOm<;A����gB�g�s����Ihp2�����{"f������̒eG��Z�'�Ǯf�G?��O��`0q@f4��+�W�/����w�H����������8� ���;���h|�	�O�Z�3��9��2G���#b��_`�J�s	�I���]DƇL�1���KH�\����&IGG�y]V�n�?k�V���}�$��z��z]AC./VcvD�O��=Z�I�0��CBW*��X0�Ӕ�]Dtp������-7Jz�𑼊+!��2���2F*㦃�� @�;���mϞ����C 2fq�D,7f���x=�܏*����ǈ�*�=ê�:Gۢ)%N˹��W��Wݗ [��=��Xw�Ed�� (��Z��PA��~e�4i O�f���<9d:YJ��q�4'�>���+Y'�M��,�{z:i�3ʗg�Ģ�2L Q������@�(�����J@Z }ݓǪ�L�z��g��JP>]m�Yfg��8�Èl!�� p��hA|�%\: ������OH� ������˗d�שn31(���=�)�N3�D�>p��*[�*�+~�MCL�,�YT�r��dBߨ����B�~}cgT7���͢�X����X��(?ڕ�N@enc��B�HQ"j�u���ݾ�3`�ʴz�}`�W�첔"F]��	�@H��,~>�$+F{ �Xsލk��C�'�	@,:h�ĉ
a �H@,֚GYd|��{�rQ��=�T?�7�.���Y��c0���&�qr�S�M��"A���=O=󬔞J)[�Y��Z�y�p>�މ�<$emll�VC��Ǯ]�k׮Fww��\"�a�S��R$�k,�~�}�����U���hFV+ga��FNh������AD`������zd��`1��A\�)���Di������#X �q���8�c��P&y�O�>�]�����0v�b0$.F�1)��0h��yX �����F;�9�`Ļ2�W���R2iW��OL	0�%4��K+0�;����:�gO����{;*��+ ��  �s�}]ʋ�Ѹ���e��9�8�}��l����;B�ғ7teie-��@D8�8!�hL�g(fـ�&��W����vD���D ֎�Wgڲ�3�㚄�gB�aS&⧝S�R]���4>C�N~@͛q w@
�n��I���K!�#k"��e)=��GFli&��w<��!������h�h�X  ��%�i|�P�J��{bN,�j���S�NE��>8���{jG�f���.놶��HhX̜>����M�U[k�h�1:d�3K�9Y�����̶����l�49���ϟ3�!h;Ɯ�޻���L4A�Ҋ�%�-�0ږ@��١ذ���q ����5��AtS{%u��U#3k1������h?>�]�Y�G;e쇙�|������W���zi�\=@�L�NPk7�\yP�W���,ZC|��f,")1R�L�J��x��;��@�2��A��+\n�;�:e: U�ޥ�$-�wCm=��/�[�<�v��m�l�	n����M	B\��R\�>��Op;����y	�U[�?v5z��	��kExGE�7oމ��)���J!�r�S3V��ů�K(�����ĕ���N��'TnV��&����&h�ͯ?���~��"l�>ONU"*�u������F�L�2a� V?���HPf�q-mY����(��2B�εh��V�J'!��L���@K��Y�rO���nA����q��V��Ly# ����U�������hֳ�OV���;:��C�YN!��*jr��K�O��>F@���q+�&ʟdil4�j���ܗF861ibB��g�t<�:ڢA���FDВ��A$_Z�6�f�xE�fXP  �����w]�������zS�<�>3�I�%����j'�FG래��6?=3S��v�T�%]g��?1�����,����N�F�#�ǘ�Wz�E7>]Ih.<��v���/~�B�,�+-�իW�@�5����bxl�k�Cg�a6B��s\2���Nt�3O=���>W!M�G���c��AXpu�4v�D����V��F��<gN�����&̼�ϟ�Ջ&������:��wmM�x�� Z$`�2�@8	����{h�R��jr�Ee�%%i]���WK��1���sk1�!���m!2����n�H�(+^��u�H��ʝ#� i�(Č�ė���.W�5���t�7�F���i���$M�U����M .��g�cZi#_�XQ���^����?�G�KY��CfY�fqVJ��4���2�����U)F��ll�޷��!h<�'���B如��m�=�ԓ�GoO��s;&����P����������,��E�g�|A��'�MC(�jp��9P��43���6��|f��iOu�ݔ� he�㍲��T왼ʞ���t���P0� b�?����NO����i��������" ʠ�g!��x,T�dzT�JcpX�3/f�Dsfd>�?Z�-�Ug[S���r��?#��|0�<~��`�-R�a	ǝ4,�;J\8��ݗ��Nz�8����cY{��Qs�H�'�0��)������/�М�F�#ҔA4{�����@�#�\�%�<���	����=��ڀ{ w�cQ�����m�~ �?�(�|�'��$��7�bA�S��㧄�A�'�&��	�-��zQ���ɚ�7�o5�I��F���;"_�z���E���eR�sه�q] ||� W"L�߹O�������C�0���.|��,�c��ДL���5����W���3�����kk�}��7ά�Y-�pF�m�o�^k�UJ��e@򀙺���Q�_�C��O������:��%HJjbY����FL,���X���һ���jk��/`��J�(��/5:Zft�1|���=>���bn�� -.������vP�X����Hqc��1�V����]p�@�� b�_� |${�j-_���� ?��e���z�O����h��W��� ;x�A߸����@�0�����K-c��C;�>�T����R�k�0��������,�1	�U�5����#t v�J����DD�]��������`�O�{Z�\�����+�� �ca��i0�'Cw�c�؅�)�V�3�A��ŭ���Ih�n-K��bu<eS�Ș�.�)��8�c�и*���$LpK��𽊨�b���@�/�J"tRE���}����s����*�>�r�w��暏��t-�i��8Փ��I�;^F&��Ⱦ:����8{�\�������S�q�)ӟ]T�.^>X� ��r���;��zQ��}�ʳ����/
�U}��Ƽ,-��%`( 
N���(e��UU�*�N�^"aH���VY��:�*�َ6Z^Vi`�=X�r��^}P	��ي6�&�����[ �6Ξ;g+ ��W����("� s�j��:�5�13�ŷI�+čO?���/�y��x�һq����
��b�E�� �J
�:E�H`!MpWL��Gu�����H�W�%�1���LƝ�٘[��V��=Q���5��_\�k{18:��bxr>V��W�Dc����lt�z<��-������XX��J
ղt�U� m�"��(Ѥ�i�ߚ������4;_��/�hkZ�CÇh�7f�伓�%������G�C5�Q>P^����h7[kk����^�&�����RN�t�]�䐅���]�(���@3g�E'wi��	�x�
o�k��23��9hA�*1���H�d<y�z��fc�[�'�E��6�io��GY���/�� �G����� � �ꚪ��C�'UG�-�N�@T��@��-l��[
�<Z>"&uD�b�yŀ��q��ngg�cD���;���;��?�a_�u��(���u!H�]�O�Y�t�A2i�P�:.ũ#Q�i�3�^|z��*�oLL��POg-��I���9AO���"���D��('D� *F�R�:S�1�X4bB�%@&�-���KZh�D��"j��~�R�Syy�$��IǕf��c ��T��J�9�⢐Ƨ�Ȼ�ځ�_ �#��	�'c�s��}��<��p�C��C�:��a���U��(	2�?{'���PO	&M�e��9ڳ����&�n;V��ho7�yf�������a`B-eu=���[_h��q�Ç,f��4v�/�޽�s�%�_ GQp��	W��\K`/�t�`p������MY)�e��>��G���͑x���_���(� (u���&�}QL̮�����v�v�㠼%�jbf�8���̊�~U4Ea���/�e!�$䴄v�%������n\;�S�E��>ѷ�x�������ڎ�����]rjW@9	ݞ?@��Ϭ���9��P�t�=<��O^���q���������]� *ּ�^��֘׸�X��X�܃"Ƙn.&��:@N����x.V��	&�:������&~B���|���#	HAy@r��P"��9�f� �F�9�� Jԋ��>/�H�ʈ�I]��R�7'U�ܒ�!y��?(e�cz�������������y����yF���Ԩ0*���Չ1x! �f�`'�~ �1a�W�% q<X	 =��uLd֢��Ix���: �I��eDހ-�@�{pG� I� ��t,.@�щ_�r0I�y�|n�<�R�U������e>��hL�d��QQ&�0lIÐ�2��#��M�%L�Ejw�:�9���=C��̼�l�s�g��p�Sv�mn$���R�Zs�ǒ�JǉS_|枟�x>{��-�9�VS��_ʩ伳gr�����;v���/볬�wE��Fv=*�>i�ҸtN�	3/P��r�$�k^(s�.N���kW���S���RG(n���y�C{k~��]i��`�ד�L���Q{BE�����=����/?T�k_�[���x�qx)�gdQ��^Q}��vF��~QM,��ލ_�������G��C�pt-�l-DICl��֎�*���i��J��a��ƨU�C�K��N��e~f��%���i��J�z� �H|�,тU�4K��ƞf��)�����~%!�>��訕���#sNXC�� ����%��_n�<s����� ��X����`p�����L�jhh����1__cPZ�O�:-˱�x�\�p!.^8z7'���>uRJ!��1%ڪ�Q�w�FN�C{[��/��==�
z<������-u��h[W��?(���.'K8)�b����꯬ՄN�N�p��J|��1=�'?���?������L���g��a����1&M#?�
�5�3 ̲4�5U��Ҁ�<���2�}��nǃ����_�������;�ܫn�k7=]���IU���N�M�h�I��F˦As����'$ZB}�5Pj%�hܚ����A��=�@�~�νx80�#����'Ιى�s^<.:���?(M����y	򺛘]4Z�A-	�/�SF�S���s<�v!�9t-e�{�&�Q� �)/6co��ˑʒnI�2��d��/���˪_.+�e墜����~�TV�����|�ym(
h_����>�{´�i_$Kb}s'���ȸ'�!���%����ɋ�11
���ϊ��S]!P\V��F
KWW�WAD!!��e>��(m���Ou�~\�v%����ӳ�Q����jU���#�ͻB������	�����؂O5V��l���~�-n���ZO���{�18�K�24�&Y�(�c�@��4�R�'� $�w3��.4mh�M`��u�w��-�V^E׀+�[��5��������'� ��1�C� �V�*��"Q:z	�8��JҖ�����_�9%�I������k��FFMeQ�h�RWO=v1�z��x`�NY��}���Zы���U�g�}V�{��Ϛ_����]ݝ�Vݑ�O=񘀽Ye�B[��b�\P��OO����%%�',h6�x�����pIaѫ>�C�v~y�,���S�{W\�P oLӞ6Mu?�n�cޢ��	���`�;���D�1N&ڀ8���N�,0����@�|-�Y�� ��ь��mm�ν����<KH�9f=�].bO�#�ɄK%�x����W����߸�`A�S6=Қ2[�ق �;1/�����e��J�=DĞ���X2��@��C#E�d -(]�1�6:�m*p��J����B�䫣N��	}�詌ui@�@���S�ʩ�{��3��y�'ZAb�$,٣UgԐ'�+K_u����Me>�W�]�|���);&�'�o�'�v�%ad-�)� @-"gR��qvVg��� i#z[Ƀ�j|40��h�|[�������x? A(>a�'��9sF �m��>�8Ɲ�6�jj_f��"�S/;�e.,����*��U�QV���֊���齹�7���FW�il%���������p���P<Z����d����:��L��'e�T5J�oԻ��0a�XG�
�Ƌ=��J�i��_��ͻ���68�8rf�b)��L"|��-�ʹ�6��{�u�����o[0&B��x�(~~4zXB{,���k�R�k:��տ�:����y�sį��"�0Ȏ�΃>���"�5�Ŏ��z�ɧ�駞��'<����~�!�ӧO{q������1?��H���~���I��H�!�X��h��ŋ����8}f��<m��i)64t������EK��u.�}m�9R|ۙ�@����s�uf����:G� �#,�B8w�3NK�����_�o^�#�K��%1���Z׋vc� 3�\ڈ�I���[{��.	���H+q�(6�օ}k�R�Dl�*�_[E����S�S�121*1�|�L�F�di�h��l��h����>�����d1.����(_J�eIx��KݣL����	��1L�ڟ����5n�,���`oDg����Oo���:^��BQ��^�䤴Q4�fq�x+�Ā���|^��ս!���1�F�����A�&g�
���L1*#ֆ+�����m(�j~��\ ��xf"��{�����?�y�0{�a�T�[����['t�4K\)���-Ԁ�m:V]`2"����y�n-��$ݹ�0>��F��.��%A<;~Z=���D'��sgN;r�wB�\#@�x �g�����|C
ˬ�mD��#1ں��K�pܺu�4����f1�VL�,��h���Ui�Dٺ�er ������+Z[{%�b��4��Ui�K1�������bf%bvE@^Pŕ�J�IY���X�R��3��d�ȡ6K������,��' �%�Dy����BJ�p�̨s$�z��	KB{@���'m���s��o��s���eR.����G_�h�(*^�CE���S.T]i�*���P_f�;�{w#f'���Χ11�wo}��Z��{ߏ7�x3>��C��@EA�z��=|�yh�Q����Y]Yr���3'����������q�ƍ�胏t�0���l�P����;��_�`!4<27e����	xP���#�G�!� ���Ս0�YX�����S�YX��j�O/ƴ�Ss�19+:��^�\��[������=���_ѹ���Eɤ���4���ш=�<x������{Q�Т�Y��w7E$�j�|�0Rn��KQ�li�)�Yzۻ����,4	
����Ȫ�Ì
����m�:���=���8�Y�S'��o���Ժ�^yR��L��4
@��݄6�-0��,�­��+i޸�Ԣe@������a�&��l="��L뒞7ԁmem�֏��8���`aɇ��*k��@�ny�����o���Z���[����E���|&�O��2�zݞi ��)/���7�J�Ny����-�-��������m_�߱�)�޾WNݱjΜ+/M��L1�k$��+߱�L�֎���oĻ\M��B����14H�a���η���{�C������ ��E`�Z}D9��7"И�����o�m{��8������g�����߉Sg.x���߈��.|M�H��	�PC�!���GAU�I�a�n>�z\���3(D`H�E!t��<���IH�h��U�v	Id������������b�#MW�Do���$�L��M�%KQ����Y�};�ăLRC!��>���>��cފ��'pѧ�;ir�aow�x�����e���j����!�Jy��-��ۊ��U	���j��_������?�����(�^����U����ɳQ^]/%l�1���7���{����֏ߎ���5nFGcei.N��g�?o����ț1=9��8w�btt����])�7����=�t<��KW�q�A��^���aRET
��}2]l�G�41�'�����.J�h��R3�M�7�W���<���}R�\�p�X�z$�2U{����Zt���~����������ik1��s�[��&k����{?��+��#�1��iI45��Z���M�7���K��JҀ$�H���-PRV��0՛����~��J�Z��"<fg:��%,ʌ����_fMUMlHC������$����lVfd�Ahnp5(���w<���0?�bDC�TC:���
Iq atr*���x88d�O@^��!�������t�d���ɉ	�S�!8�\*D��y�
�ӑ:Lݘ�P�2},;���f� ����g~Rb������e�<�W{1e~���>.>�����_�x��G\hۣc���ƭ��(��Sf��8�;���ج_W2������G�cX�����U쏳���Jc2�����w�̈́�]��87n\7�^�"�De�C��h����]�4л-:s�l�0��
zU�Vʺ����j�w��W�+��Y��G��#��h$�����Dɠ�0�e$���<"Ql^�Lm
���LY�3L{&nI4D)"���DF�:�ͣd���W���?�,���+oy-��%�Z�����]���I&�z�*	W"}�7�e�˒ �Ѓ�J����](^mei4�WGk}� ��_�U�G{s��/��ŋ����k����2뛱V�e-�k��8%�C�������Z��=/� ���q���-�4<wdAv�]}�NFUM���o޸��/ǡ�c����|��{�ЉtJ��^�*m��6%pwԦ{�Wa�AqylJo(ɕhB����E�,���yF{{��Pڣ��))W�[¥
�_��4�T�}YhHP�"ұzP���/^�_U������_�O�A�3��x]L��=��v��ʿ\r��L��V���`t�H�w�4�ei���N����wi��U�b]���E�hq��2��0ퟏ���VS���ai���cv-���6_%����H�<䌐�/L_�آ�4XdA���G�p���B�,t�P�Z@�&/M��QOђbZ��$��������T����[�Eڨ�S� Rʎu�b��Hn@��a 6Z	ב�յ��W�C��  �y�KX�V�F=䃚vK)�NƷ�;�rLf"d����C��L�O����W�I���v��:�4��O�}���<%�֞gE{$ދ�T�6a��v. ���\�ڥHR��'�X��\��"������gxQ;��=Y>jf�r�ǇX� 4��D~̩ �3�ט����Nk�R��+A�	<�|UV���6{>P��,�}������p�R������x�����c���K���x��x�o�w����o<��x��1�H/���!><Lױ��޺}W喕���o%�tt
����>���q��
�$	�ߔ�%��ڃ^��B���SO"��'RI���/S"R��&}$
�[:ǂM�v��[J��;�������o�k��  s�4*�����T����O�#/��'4�TQA�f���hi��cD.�)�̹J���&�2�Z�@�Ҏ���A�$�U��~1+}sL7d�'�{/J�o�E�*T+��v:���n�H6��<ӿY<��M�7S��30s�ؙ��C�z~R�H�P�.J���� �����&&+�F2�xUMLQ�
Mԫ�K>T��$?&��ʀ�����P�R:�x����;m�׎m�E>��
�l�+%�r��f�-�"`i_|� <��6sG���@ b�	�$|��/��=�l<����駟�g�}��X�����=��ܳ^ ��	��9�,�g�O�]&��i#��ȣl<�ꊉ~��>t�+�O������/�-��ڡD`R"�,��^��Px�~�̹����G����
���u���E.�*~a�����X^\�O��ga��xguEZ�����kW�}"}V�;0�V�N�>)��ok�n��I�H�Nz��E ��EN�{�W"� \F,�q��ո�����O�O>%a��]���&�ź��R�m�k�� W��@�s|��u�?ˁL�����t�a��GC���j��@����ϳ$�y(�1}�Gͩ>�=�F���l3�6�����
S���(��'�0dk�4��ݣg=IK< =�ݬUFa1qL�!�x��?�g����D�O�E�4��m�!Њ�)z��	��f�044�e�F�JC�`�BASRB2�S����3՘=���*�x���1T	� q�)��A*� �okn
�ʅ��5���{��0��`Q��3p�i�h$�fFU^ ���@�b ��n������s�F_)!����>�w�yG�p�&	�4�C\=��10�G0�H�����DV�d��.�3A�������µc�}�K�(�raq��Wo���qsݵ����O ź������l`i8�o�+2 F��̆f� �Л���b�Ϟ9�g���w��Ÿp��#9z{{�s���8%Ͱ[����q�ҕ�z�Z4��p�?���۷n�ϟ;�`��YX��+���Ĉ�,���0&uC@���c�� 8_��N�{��. u�7j����e�f�|D�,���0� 	��a�D���.�J�zd���a���cG����ΜY�XB/�'��u�ӌO�^��pUKeQ:V*���e>e���L��+��+ /��k�ai��B��Q>Vg�a�D�N��E��٦��hn����V/��ZNDư&>��}r#>�~�.��W���"/m>44�=�|455���J�TAŢ�|�gbr*>��z�V����.�nݹ�/s�<uR�oe��O���ծXod�Q=U�Fcq��9��u��Lm�>��(���;A	O�a������%��͍Ŵ���(���Rx���/����qyU�W�\]aQ,�ߡP�"	&¤A��ed��+���B�� >V@H6����&�j/x���~O -�B�ƒ�c���[���.�;� ���~:��R z4���
5� ^���q�� ���+M!E&��!R~�vX�_�̼=����A�Jc�Mƫo��çf�e�Ul���	����tv� N�I۩���ѐLܣ�K�+vaH�63I�����kǷ������ڔg��/����n	6q�4C�qM`�ꉬ�O�%�U?ݹs�q���D�����D��o��J�~.��.
���,��򔀜����,d7::�f��,�� ���b�L�.��Ν�ʿ�B������	��E���zeqB WI��kj��� 0 �<��1@���J�ط�{`r��/� }��w|��<���+�^s����Fj���d�&e�ߣ?�3�ƨ��n��}�ĵ}�]�ڒ��qi��2(O%h�z�~P�]��WbzG^�	����!����y���S�4��\�o�V�_/�#`���v�,N���Ø�K3��>���7,���'-��>�w���>���N�Uc����|��o~K�Zm��8�K��f��
��Fƨ�d\���Q�����7>u+�&���{�Z��&P^�X��SR��6`p�L� �Y2/��nW\BD=�Xz�<���B�3/�� �Iu�3 ���=�f�ڲ�T���?�O�FiEm,�7������cp�P :���)F��2:Ѓi*�J�~Z��B�HT(�?�R�6щqA઼Z��� ~
���q�P�4�z1���0��i$Lխ�u�� �k?�+i����tB�xJ�4&�0�?����\|�;"���i��"��

KD�h�Ф�D�HC��u>3��~`�!��6��8Z��.�q��܈7��q!���Ǻ�ۗ�����e����ꑄX3�^:�G�^�tx��e��d�B�Ⱖ
�g�C�zִ��ig����n���ƭ�7bzj�~h4U/ ��Y	
�c�D�<z4�5C���4V%��>0��;%����<�2J�/��(&WB��Ǽ�2A�J9��*���Y���7�������i�N)=�3bx�"}�!��W�S�am
���?���>-�f�6ޚ
��5���|�:�)�z��I <���ȵQ���DX�**�v^(�+BKW>�u�/����Uлj���$z�
� Δ۠�sa�r��Tt�K�1��V<zp;&G���ø{疿��b� �Q��Ѕe�>08�eh�z�c�t���=L�
!��|yu�+p��/x�[�0�ﬔS�:h���3�\�O>�D\�x�A+�&c|��beˀ�D��n��'{e��!�Y/�q�̩8��'z���x,���V��4����0Q��d��5�7B�C��G����9&�������������Fi��ŷ��'T�4��t�/�9�g�`E?V�����m
B��, �A	��y�	M�nu;Đ�$[��Ң>,���������8hH�v%�;�H7EC(����X)��g�8p�f&H@X��0����Ť3s�z嵷L0�����Qڱ^r&$z7�t4K��a ���P,3�D�n����5$Q��y�:0|�-{��nz_��_��U��������`��g�y�!�\G�D�-��(�Ey�
�����0,1���a��u��ƥ��=��P>��3��Do\�xѦ?!��I����%�@���H�Q=D��-�qC����$ �BQ`lˠ�t���X҆a@�@+n��R�/�K{1��*֞	CO�g(E�X������=ě�H.h�ס�(r�#��
=�{�B|��Ti`�D�2��4X+�D�*��_VU��@�址:�>̯� {�D|��F(Wr��r<J5��E:�{[+�P6C�
�1!��JI!(�������;y���÷(��z���"Q|	"A���v�@����Cߩ3�\pG�Y��K2`�h:�����p�8��7��o<�L\�t!�z�<���b��_���z+�eq��,:t��@���p�E|���8'�g�P>��XZ`��$��c�g���VQYnj�����������XLL	�+��oG�*z��Y�iz�̟Je>'�qU��3�yꉨQ&�p���_zI�X)��i<3	����S! �lŢG��"L��z�#�RHg��M��ѐ���3##�$������=F��� �g��Й5c *��o)�h��3�̌��,���F�$��������4��:���W��H�4Ȳ�ĔY�))�4L��� s�1<4|�
��D�?��{m�Ar��5`by�p��o��G>{�'n�3����y`�� *ij'���ڡ�p;��/>/(��櫫oT��$gJ>[\';����t��
�#| �Q����^�'�氿6�:��������� !�f%���i�Ġ4�������fb���3g�\��� f� ��,�NV�!�x�c�w����f���u��u[�ڻ��qܧt((�9��,��Q�p��B��.�E�C��X1"흟�p2��u|�W��-ހ���)Z8��7�-�iU#%2E��WP���oU)�-u�70�!�y?�u�E.XT`'�6�"=��1R&K���<:Z꣯�M�q{tu���;:���7�:����O�'=v��ݣ�m�EC��{�q)��~?�G���]Ұ{�i����p:N��.���Iy�:`��c�eyn�CF���͗���Uy�l}mKY�m`%q��_��嘚�W����\����p�rnv*v�֣��9Nt3P���-�Y���a"�����4�ky��t�
�V�[_%��G�Q�V�KsBc�+Rh�W�t��/T��W����g�^z� ��ʂ�5��o�e�*|<�į����V�bvV�:�JC�i5;Ig�������D0��B��	��DHˋ�j�����r��F<7�B��4q�h ��0��0��=�Bb3�MLuI,��Y����[o��x}�;d�Z���Ԩ� �L��vH���V���\�3��2�"0L܉�%C�	��Ù엏|�s[~�K.}fKy�y��nBځ6��:F�Ư�B{a�m�%6m���舩^XX�����B� �\l6�	�䳉| �DOW�ʷ9�Ĵ����|��K��<,�2 ���WXkxE�>���˙3g%D�)��&���|���'�:s�8r��Ǿ�g�k�Qo�ғ�79֝nߖ݋FD'�sNH���/�특�n3ve�S�:\7XI���䙱$e�wi�la��h)++���W�%\<��&�4��a0+�+��̘˞��w��ζ���䍦�b���Di�W������M��^�/}kG�A�4����8�W�������:��)�OWO_�8y:�{OJ�w3X2�oE��xW�^��q#Y�&:�V_7�"@:���3Z�ڽ:l�����4�0�^�����]����/�^e�ٟ�I����V��:ڣEC���Swn?��wnzr!�2�|�B\8���������{Q(li�E�	�?�z�����G����\JO=yF�`�3�We�0`̤>�+��\��������D���,�"�-��&V����_{;�}�k�׮\�˗OD]���2Y���$!�ʸL��EiL��w���0Μ=%1ea���"Y�Ω��nÌ|~M]j�O�&��9��fy_4�}��(�k�7�LJP1a�5s�K����X/ͯ��M�E�:/%�����PM��5I;c�g���R�'s
��6�ν���o��n<�9"Dʢ�Se�{GEI,���<*F�4�����`���@�C� #�G |&�%B&/��<C���73�6?�5������}>�U7��jd�� �v�!^������0p��8���������ͧO�a��� ��2kD�<Ļ��  R��`y���y1���7��?���?3���^���{��{��Uk�,̀�[A���A�
@��� ��&�O�An��ƪ/�|u�6���N��m>O��>,��SYly�:~i��)µ�#@f�Ju��3�W���~y�[�"  jBg��ay �LZ�W��_M�^��>SP>\�ź@�Bq��= �P 2��S���g����i<�X��"�_:B�*-:�bvlI�I0m��׊p�/���@d���ʺ�%�4�����^���Y	��Nʑ�P�V]p�h�87=���<�41%t�oU����|E��{�ܽ�o;�w���xL@���7��^�;����+֧���˗��n=�����Sj�L�Oo|�I|���Q+��'AD����H|"z������f�����������>Lhd�@����T���?��/?�ƏFêx�P�6W��2OZ�T�o����2A�`���
�Η��wr[[�bG�����'e��<����T)���X q�,���s�7Չ�<���DxLc�{q��y��YW�h;���ӈ����~Y����y�M��X&bG�?L�@�N�}��ü>��Ӹ�`PޚX�]Q��$x�&*�F���3��#�_���sg�Hp6ƌ�/5����$���}z�˘8���S���՛�
��6��Sr�ٶ,��<���:f�Z��.j#���, ��M�뢁��_�t��DoiJ<?Q8X��D4D7J�+��)��.nť��X0��?���1���� >����_J�@�ȴG�gY@��e>v�1	�v�̞�#Yߤ������%�XE�(td�U���ф��h3�(�w��f�L��s����^u�FwĚ��a�OJ,%�:�a���12V��oj/�G9�>��Aн����f��Xl�k�pA��S��òX�X���-0�~O�~��+?J���"�*q%��|9O9yM��PgTI�(�ǅ�3��1��A<���O.&\�5����H�{�B�������S�䝖���@���w�߳B�����~(O�1M $@ۿ� ����ɾcM��s�<�O�9�P��؈�h��?{���cB�������D�����y������,�����ht2u�щ8b�9�ɫ�]u��,,�/.�z��C�i	�%H婦L�n�RG��T|[t>�
�#�vv��"	'�0̒E�*�uғ\�(1q�)}'z������I�H�x��n�MY�FJ���-b%o�Kا�� ��q�@S���m��F3��BZ����ō�uw0�|����+oǏ^{7^����������yg@�?�>����'7��;\���;��(�|�x���q�8���b&;�A��������8�yt�_�����1cz�R2����}�� n��َ�罹쉟��ҧ
egҹ/T�klG�L���ϱ�٘��o��'�x�1=��*�%��g�E���7�0�O0�_}�����o�~Z�lGhc��0h6>6�� =֠wQ2�h�h�	�Tbxi�^J���=^��ɍ��j!�	Y����;v^���Y���%��ܓ��i����Nn"D��lN���tX��F{ַ�����O+X[������ �-M�B	�UF��d�Kuǅ�,Q��p;ح��v�ו`N�֪/̓�-�ǡ��n��y�\= <3὚�;��ܦ�C�x�O�����r������'g|RZ��\L�1�Nc��q+,�F$���1���C��w���F5yh��S����R��H9@�Q�#�K4�2���rI(*O,	x$�P�s����ԅ�`�q�a|R	ZŻ�&O�fG�0WY��E𶵷K	�$�,���-��0W�	�o�
���<�{�=��'<�1̓I.x���#1�:}�h������E�4c���Y}*�@4t�H����Mho��z���" �V�PJ@�< �_d3�8�Bf��DQYMl�������7��[�16)K`z9�=� � ����_�q�����ޏ�����'2�Gcn1�_���z�<����t�����?;��gw�Gݡ$Lz%��kNٳ_�q��ίL�=̟���w�ܷT�ϖI������b�q���9�	&O���sФ�~�Y��!�ϓZ��s{+!(������:"����7��_�_��7��ǯْ����z�G*�;B�r%M�c4c@�rV����姶�ߠ/e	�7�k��0`ȋ�Xfɯ%EIψ�_�ʪ��#�,�^�z� �4��/����	=fN�o�:}�\F�N4KM=�E �`�b�_��Ю�M �MUU�W�$p��j�Ǚl/.M�Հ�O'3b�zȗRH�}�)�]}��9>��k�2	�I_#�>X,Y����uLD�I�ˀ,w�6Q�z�� *�'*�������"��K/�s�=�/r�&r�E�A\R��T��,"�O(0�����m�o��C��V;	�����\�^ٴZ���e��E��3�y�ځ�BC	tX_WBb�?<��1�k+��3��%Fؘ����. ,�V-{A�<E@*T�
Z$)/��t��`���w�"Y�@ӗ��s �H@��;���k�J��~�v���q����|��	�0�iN#ChN*�j��?'��3T�5�d+�DyUm�6�DYU�L�i�QVY��.DQZY쯽�n�������{qWfڽ��`q���U/�����F-���.���h��/::���Ք�����̑��H��>�%m�����'&��s���k%�??�_~g���3$o�@j;<�+:�vh�M[�one�uE��@�%�N�l����g ����0q�q� `�@��I��Y�Y	ai^Lz�]ѯ�GӇ��R����9�L���3h�e%0�
��]R$���*{�ճ�	�|��#|�����Z3W+�P
N�(?癥�V���Y,+�	K��-K����ER��R�������M�8
dS�Ue���B�8JtRk����q�O�e*_I)�Z�y�XkIy�)-�E��V(��)k?7�����+�y�Z���	�p, �ǞaK_I ��'M%�8���ay�?>��7P��V�<���pL�2{Ot{�>U�"Y|�e��$dk�mUʷ�n-&~�hi�Sg�G�IY��.Ƶǟ��Ξ`=���cn~=N�:�uOSs��?��v;{R�h�!n�>�Y�e�dɼ���Rb||]��q����&������B ��	]u�,&�,n0"��DcKW��p5z��Em}��K�T�+��ҩΫ���f����x���L�d�I_\ތ��#���7�7?�O�ߋ;����+Z]Ӡ�I\��`�L���$E�a/��a�=Sf�0ֻ)��Jsk�L������TП>9�x��x����+ODCk���������=jZ���I�S��/�&T$�pa�]Zoܬj���3�D9ъ���%P���7=�z���Ov>�����61�ӿ��o����%�?��W�~�s}k��/mb3)��l���btd������v�'(�>3Cq < {�!�Y��������?��x��W������3 �	Z�q(&����f����ߘ���2kY[^;��~���̏k����w��cW�s��������d�����[��4p�i{cYZ�rl�-���R)/R.%=�����>�������M�+��c!����u�?S���Tg��w�u�5V�Le"yݬ��Ǧޱ��{�U����2�Ih $�H*j:b��H�/�g�	m��y�1BK�=�������$4g�1g��^ ��p��-�%}`)}�!�`,s���@#R���gaa�A*�Q����Pʎ>��fܼ�PXq�����������G��/}[�^�U~��?���)�M-��_������?�}�de�-�����@D#ʒؓ��7R
$`
�@/�n�)�7�=����XXQYԞ�+�``�3�����ED(� ��^���(�n�2�M�-���h�2�ťOU^Tf�����a�#��X����Y�Ǣ �[�V��l� ����]1�L>=OT���"��E�����@��_ڔoCfо�!��у��8)]"J�.Y����skN�1�hH��2���@��d��*��Sj�!$x�R~���V�/nb��K��?1q�S���7�<��\;�_�5�����t�{����z�0;���?eKw���Hߟ\(#4󅯘��R����Z=|��T��Pܸq+f����Ɩ2����M��,�0O��LdfM65H�ѻ�d50��g����Y�Yt&�cEFB�az����IT������\1���Bi~|Ս�=pһ�bi� +�|���am�r!
�ـ'gm V�d����+{�gO��,@I�@CK��%���ꅻ'�O��Ț�=ybX:n���	�}�����&���wX;�f�i^(�e}&���E�zZ��'%/�K��.����F�<�'���Ċ���X���`[�%�nz�%F$wb�Ε"��-{t�(-���Ο�^�F\�r1N�>�=�?�y��'.^�L s�D�(�Ѐ���u	]i�D1nA$!���H˛o�_�a�ȿ��(����M4��޸�E!g�%�
�����֕��,ϤE��f�a��8PV������/�̀<nLd�.W�����T�_T�`�T���3^C�3f������!Fy�aQ���fg���gE�ghX�dވ�*�cFL�Ꙕ"rlQ�@�Q|��3H����ܹ�^@����E!�}YJ��B�3G~K������AI_im��eNX��'���J�#v`v&t�v҉l��<�N��/����~iED} �|4fJ�)S�YC�:b^RN(�>L��ϱ��9J������������e�H�>{�7��mr��촇�V���H�!��|�_흻��^��:q5:W)eC	 ��CO�{B9	�#��UZ��H�B��4\9���8;?'�gY���@��0Y,�55�&*�={6ZdU�t�M����|D��4�F�E����s֛G{,*�v�V���.	mf������+\(�g�ƛ(5QG�4��Ps�{ \���P�E׼�F��5�h�%ʗT*�� �=���fY�m�-�d�;(/�՞�%����ɞ����yʆ ����!U>�K}ɞ>G��e�oJI��YgeN��y�QO�
!$�^�7Vԯ�`�T���Tx�,kёZI B�Є�����N����ֶ�x����/�'O��֖FG*��%q����/
�Y�,s%U8G,I�⡘��7�����la���{��ӛ���K�k���#�J�J4"��'Rbnܾ�5��
cEM�^��5�}���ά�m	��)���.��b>�my/"�*�4�ѩ�(�j���Rr�q�|���L�v| ����qeюY��G(���u�C�2�>�(���| �L��NW��{!85�.�����}i0�ĬW��ԱzN�g�\����v��Z��r������8$D��E$����x�I��E(�D��ϯ�<'�3��y��T�j����	�UV\G�P~�T:�x䓎���F�)��٨Sv���>[���e��) �o����3:&>��J%P!���6|	�-1�ÁA�J�}��j����o��E(��~[�KbKiwk�_��e�Φ&�����  ��h�J�!�lE�a�ĉ����56�Z��K!Z#��~��CM����S����4~���`�{ WV�L��Ų%P�Ͳ�r���B�7|/�lcm%6U�\2\�Xs���y��@b��6<P�@o�*b.
��lZ=G�,�F9p�x]#�q8O�M�Qk��38lL�����S��.c����'^&Z0Y	�e�=Z8|��UVΑ?}H�95��L�q��v�>YT}�$(��to��qq�C��?y�1
��w�N��g�������hif�=�-+�'$dˢ��g�����A�E��F1��[ʓ�b�����]�H�C�E,^W)���[�1>5�F������#=��vS=KD�m��ϾN��:t�ӛ融���$��F�ɻE具iucAX^�6~�����o����]cm�(�Ɔb~nZ �x�u1��@��y�*&6�c�"5 ��Y*-��L�$�SSZ4cJ�eL�-C����.L-�証�  BI���ګ�2�t�:�
_n"=m�@#�y��4��)`����z�T�,��b�p��PF� x4�?�!��e��K�b�M��Z���7�7��o�9���|�a|�/�<F�GLp� �QٽvJ� ��I����:z�Wn<�u6����朔���1��<�������h~h�<��:hj�\0��eȄ����J�j��}N���ֶ����ŏ^{Ӛym}����X��ș5�
� >3'+���m$W����<����ԺT>x���hh,�{���Z����1��FYbW��(z��w��}g�����{�6ju]k�5wFeM�-��M��H�倉p�(/���%YW��'�B0G�]h� T����#����Z���g��6�Ц���1~q"u��!�z��k[|��<<T����M�-G����hk�Q��;�k?�^�bM�Np�a��oS �/[��`����Tv\x9m�¤鳎Mi�n���	Sci~�k��	�g� ��y�:�.�3�����S}$B���>�*�T��x��'�٧��
)}�Q��?����$��٢g3�� �D��B:��ܻ ����Y��$��ָ���+�\�����IM�>(��WQ&�0!|�q����q�� �IvD���e��=��&R�Ƭ.Z���o�������O�GuCw�.nH�G���צּQ�1�( #ߎ���)���ĬrL���D sb�2�ʘ�GЈk�{eq.f��.����MZ���������$@�����HODQ�r��\�1���QUS�|%��J��T,�3J�YN&�c�E@x��Z�{4%f��8 G?��G���	5��)��`oC�l�S�?���/���g㺀��W~�:�i�3l��p�8LY@0)?��w�n�?e�P_c�:w�Jk�_c;�4�q��_���m�_�Iԕ,.�V�3����������]ϸ}�o��(U5���"��f2�P+�}S��Z��Q��R��ʠj�:Q4[�����W�~;a��,Ld�e�3Ygr~-�:N��.�����,�������q��ei[+����������ʨol�چf373F�o����[�;�>��ى�>U`���Ћ�����?��6���ad�I���U��aA.(8h�������+��lI�H� ]2(��ӎ�=y�M���|3=g��.i�X�ʒ��pP�p��J�G���a1�fAP,����+���s���Y�,bmy1��Ŝڳ� �Ghx8+�6����ʨ�Po��n&PR�#��?�O�~�ǿ�;^C�����}���w��x����
5�4���1
ZB�F�Ϣ�s�Xˉ�445Ǝ�vPK�
-zX^�2��̯H��5^1@pg%-���>�EN�'0��W���V$hS{F�./�\�:W�[O'ga%O��T�-�9n����{b�4�) EpL��et� 	M���̌a�����7�f!��J
e&ω��J�
pg�
wO�,�#dL\�sh2MD��Ɉ����1 ��D¥��VTK+1:1���`�F���2��,�� 0y�/�{w���P��9H��X�њ�$.��5dD��E��W��Kq�������5?K�J�Rg����� ��<b�8�+{m��?qˈ���ʯ�.��K���X	�����ǝ�	���G��E�j'�v�] ��=�^?�?���j����mRW\k�Zd��ƚ 7�������c8�*D��e�b�5��O��7�����zĺ+e^/G]�	�G�p3.�J�����q��y/���>������r�yu�-�\˦5�V����_t�ٿM;�� =m����M���0���T�����4օ�[RY�6�<=����On�|ԫڲߺ˯��Ƿ�<�(1�%�W�P�8ͷ|=C E�3��@�z]�B�R\������v|2�����3��u�j�G�LN������?Q�$ 	���%�0�������q[ʮ�^�se3-���~���d��TV�_���������,ţôR%E����g��7Kǒћ7�cG�cb͢zY��z^�-��n����r�w������AaW�#7$؊Y�U�U<�b{+�
w���W���5@9Bq@��U�	�N�����V4uj�؎�����b���2�*+S�wf�$�0�����z1�s�h���	`�����.{^�0���O�L��N��O>�_�Ο������=��Nx-�|��sJ��,yz���8%	Z�(��o�QJ�!1p[�F���$�2���O��$)����<�/��_�O�����8qB�S_����&���H��Q��.,����YErrrB�1(�o��d0 e���-�'�0-Oʷt�'n����63�ϰ��)����5��c.�����B������z������V�I3�CC�%|��Є������|��ʙh��m����,y���}}Q'sum�~���U�).a��i��;�v���7Q����m[����Dt�@���R�<xt���Ϛa]x�!'�Cc�\3]���B ]y��1ݐ�A�l������k"�#D�qJ�������$)]�߸��c�y��u<����)�gߢL,����ŋ5���yL�o���?ՙ�%π=��z#>u��z��u	��֖�Q��r�鈗�R��m�%o�|�<�� #����කf��G�-��pDπY�����Ʃ��^�����}'z�G����uu|J�TtY*Za��MJ���+(;�E Z�m%T�	F�p��R��h!�h�c�z��Q�z���݂���J�����P$km���Հi�&���46K��y�H@�'���WU�� �*�:O������-���ĵ����O���m���.ueeY44�G�L�sgN�C}ه�����^oog�u�X����i5��O�(�ɭ=AǣL�QT�@��H�n���Z�"'�O�)�!ڧ7p��!�E[��E-�r�����Q�<�$�O�48)/���ޓ6������s�T��i��?S�ϗ��槇R_p�Im�+�>�e�r��s�=�=	����!l�K2KӶ;O�@?S�,au�6��jE�D!� ���U��{�@~��)�u�X���]\U�5�}���6���������a�+>�1'��j`��ą3�?/.̉�q�;*p�����m��@)Q���ς��f��*8�x���i}�[���r��>���ߩ͏�1?��9h��|o�	���wu?0�'�6_LMw�Oy����eS[P>1�xrW�����Xf�غy�
�o�$",�!�q��u�\/��P�%�3�F�WU ��d��x�̉�+m���~PP��Ų55U(�Ix�D1?A�ްf��˕�1��ZY�����t��h�w[��(�x 8+�S�O�hi�J%�h>�V�q�^V�M����Lj.�� �C��w�c7���?�8JtP��1�/_!��PR�@`ORAq��IRU��\g��|ݧ��@�j�P#2 i(�X_[����^+&�������2����2�d*/�l^Z��M���Л�ɷ�8K��Ҭ�byI�(-/-x�;��`:3Dǚ������y"r���m�ƀ�Q�"&f�� �R�t�d��i�l�Z����>�e�|�W����!���lz����G�p��?ٙ��*�G�qjdC{�0�?\��s���FhD�2K1�C4B�������!�X���/��R<��s���l���Y �E�~SS��et�`��TP�'���q 	��i�!�|�	�>@]!аf���z��< Ē�����yl�M��]�;�����V_�;my�)�;?�oI���?�:\x���IP�
�u�����[�o3qP��A����p;UV
|�<ʀW{�Ʋ�yq~*Vd)��-�zZ�u�$�pM�>��~��O�̀hZ� ~�Ri淅�*�V�>p�)�%	:abuf,��Yဖ���) ���8)밪Rt&=��߷�� u�O�x�Hd�6��*�����dT�F�U��}ƞv���'Y_����(�]�n���Y{jǽY�Ж�\*�P��V���$x����b���:%:��?������h�N�FEMC�5C����8�BJDA�Ѡ���ra�e��7�
��-����U8�8TCl�z�`uE���������bHyK��+ʓ�� 4'��3.���R���;�������� � �4<b��4$t�r5>�btF�w�$A�9�>w�%�l�A�� ���C#�=�-�9s���Vi�h��z�v1m���!��Vk���Y�����19C���j�x�g�T�\���Ԫ�������_�L����9� =LH�I\=���X����Gv�0A�+R
 Ѽh�Ɉ׿v�J476���o!//�Y�� �z�����w�Ň}���Z|r�S��f�7����f\�x5.^�$ .��#�/_��/\��VY�|�>{Ze�y��
q��K-�	55����AC">��I��&��@��t��[%�'e݈���
�8wa�-c ΁ �b���1����s~��������>&L�{�s֩�U�K7�Z6,��`m����v	�&[KX��S
_���=�������pb�#xހ��+^Jcf�A����U¤,��ؽ�<xvO� 4�_W�
D9J��/�1V�ױΫ_/_��r�Bǰ�V�e̘Զ��%�V��#��(z��Ч��F	�L(�#׳��(om�+���ǓqG{>�Ch2�P��s�h�r����V�ZY*<���/?z4#3QRUk�VGl0Z�ѕ<5�_��/��i2W��n����&�nZ��f
������s��Dtw��`ei�b��^#���1���.IS�*�"���U/����i�A�>~=���C��Y�t$�p���NI�f�C�?�ݜ�!���;e�!t�S;��
uogG���{���gCS�����C@�.��3�1[���TDZ�p�.١�����f�'7������и�<E�~x\������7�H �aK�g���
�WUTz�f���ٞ��{i^\0|��u�o��&1˒�p��<S��������֮���p�?j�j,�6��o��$D�4�+2eRZE���N�΍x�7}���{%-��Mc�m�iFЉ���t@�giw�}��W�8t�A9;ϖ�CJG.��\���d����ӖΧ��f��K�E��BB����|[;��)�R*JaEO@����{a9 ]���i�9����h�v⽴_J�����3K���oiG�"�������e���)C�X�RVq�./�	�'czj&��c~v>��}7>�ו��9'z���p]H|��9��h,J� L����k<P���m-���T��߲@�ڨ��ZV��J�Wɤ2�Oe���F#<<K�*�u�.�����G�����| �Ά��dP��q�D�Uk��	�c�̴=I)@��v­ �V���1z�ۣG������ ���fh�U	aV&�����42LD|wh.tk��e+ֿFb��<�0����#�>�C*RV@�r�?&Ƃ�(�	�M������J���S��eFR���fwJ[9��J	��F�UY���5~�Ĭܢ��?���/�F/'u���N?}�^�>���?�/��՗��^Ͱ���_?�����Be�G$?��ښ�N���	
�����51��u���@�g��~;�::��]�}�˘�����L���KHXȌ�������;�E%܊�s�������a\L�B�L��k�C1A��i3~�{y�I�Lk�>G�dm̽�srr�/�{��% ���}��T��S:~|�����'��sI8d�G3���I�3a���2�nL�#���4f/����ܭ����=<�V/e1�I�1��Ҟ���suL;'W�}��iR�=����4h�h��-TWU��,G����G�����ݻw���q�歸{����E��G��}ƻi�n�S�M�q�To�?{J����DW���о�a9��=�m���"<m���&	
���v�����Z�<x�c��+-�Nzm���OG^y����Ƿ���;�V1y�ti����`JBK�R\L�f�)2Tih�B������3#�WVW��g����<02��I%a���_��0����D��Ս�;��Š��R�~,Ȥ�ّ�W�ϗȅ`1�1{�Ŵ��Rҍ�jjH��.I��\F���0mh�N��J��������~�����~'�\��?�(^������6Y����#���1�3D� R+�]��;��:���3���G�զz俸#o����ݕ�� �+}o�P�������'���o�3O?|,�?z��Lq'�����Sz�$E����_��wE�Ub�O��S�=v9��۷Σ��%���kOēO>���_�7�:��:��_�Ʀ�x�w�O��O��۵�@�ʎU��b�����۔&����f�Ŗ�$������n���EǾ;k���:Ad
ֹݗ\��2�ÝAyܶ�FF�d۱�����p�\~�?s�8y�J<G"�շ�Ǜ�哾�G�sav�g����(߳��)���Z�G��w1ș��z»)~�>��UV	�f �O�VVT�b+�r���3�Ѯ����cХʎk
�F 0F����b��um��x��p�5�:�:�������L��ĭ�M�܎�CVA�Q��0z�JοDC���b�8�X蒶b�.�3���MM�J�!,_�Nq`ID��U�?�^}��N�Dy��E�BEhL�B��b5(	߽']I˯Pc��.�-�����>N��+����sg�ʅ���kIE�+�|��W��:;d�0�#y=3sJ���fʮ
�|V�f
������[#���V�"��>��
)}�BO��rD����F�ԡ�C�ڒϥ!W�QΠ �a�m>�.m+IKH�5~IdB��v&�[��'�?M��{cC&�{L2l���7���m���lG���.{�>�����˘���+ �vqt���L��Up��?�����+I0Q>0�5K=�'��q�>u�t��H���o���3��|��/z��;wA�Wo����k𗎈>c�Ё���l�dg���{�14|�X@�2/	��c��y��M�Su�.z+Y�̀ ��i@�sѲ����.в~�4�v�)�g�"8>s�I��}�\���A�%ƽ�2J[���}��~���U,,k�ʃ�kx��+7-p���鴄7CyS�t���90�B�p.N�6�#���Ա��'W\7v�"��{R�D*�#�w(�h�>��r��)u?�Op�O�1�N������w�tI�ة�'�瞓�p-�1��&�����ۺ��h�r�"@f,��^������Ze�=�iR�k�u,嚥�����T�-�,�6i��-��ծw���k|?�qN�
k@����o|2|����;�����/n�`�P�����(�O��31�_�/��G�2�ՃPoߔ*Ц�44X��R ���3�@H��Ҕr�1��=� �O��;��L�l�âv����֖Wd2.,�<�p0L%~z�O扸X������,�[ �B/f�s�=�ph�&l�'��L�xf0�&�R~i`(�c�Ǔ��_��_�g*�߽�?��@�5>J�Y��3��#T�M/�Bp����_���Ɏ\�|���$X~����o_v��}���e戬�V�ꁎ`@�����?��3��ODm]C|�?�7�z�W�  ^X{�������1���7��>��ܹ�2������YP�I;�%��WTTGGg�5͛��������3�/Ʒ��m��_=�����~i��GР���[�zB���Rt����@��;՛�|u�=� ���}�h0����EC�oBS�9Ө�ݟ,�������<}f��ޥsh�,�BT��r�d`��0N�x"O����+��km����r*Q'Υ�b	�G=v����7˵�2)_�*g�b��ާ+N�[�P�0I�G�����(�M�MQ#-�e���T-�x�2a�0����cF��~���'�u����?瓉]|������]�(��4A()"+���hQcsL��_no�	���٧�EԌ-Ւ�����w�D�[�L�S��]�j��_�g��?��?xyxd<Ʀf����.B�И����FMe��J�Ϟ�ī����;�'{:��^R����n1dgt��(U�x�.KHg� O%��Z��Ib��&n"��qL��R1L9�唉T�c�E
��y�cg�tD���9��z�X-		!�pϠ�ўt��[0q��(i�:��&J��D��҉���Bێ��/�07�/<�	����7��L�sV�xG�߬����_���eӖ���������,�j�����;��S��AFhj��<m�e���n�~�?���mH��B;�*Sֆ���ӧN�y��A��� M@
�`2V��	coo����x|������r�Q(�Ï���"���n�>�B�#��#04H���Y��3XG� Bą#Z�Ȗ��W�kh�uR�'��D����9�E	3��1$�e�b܃U_;�/=�9@��F{�Uh�Z��	��w݉?���_V긄���P�����4������R�Q��?����� �!��>�\�e���J�Ke���`=��h��jS�u0�˚a�c�R,Y|���a��,BnK���ڪ����%4�p�}s/m�0@	����/�v4
�v89T{,%=U������9�C�v�!�Kv����q�㫛�{���C���k^e:����̏o���ƻ��oFUc{̯�r�4R��Lq��ɤ�m�����^k�|ͧ�T���G�aR��K��:���)	4S�����#'�4�A�?��/idH�:��!�IҒ�Y4}P	�ZX\���78gff�i5�]Y	|��ע��=��f(��p�8�j�S|���*��� v���{�k���j��ߋ?����<<�Bs벨�"�ˋ�e�ML���Q��O���������_�?�ܗm_u�_�i�ɚ6��a3��퍏�w���|�xJ���9���?�7��4�Ei�D�H��?��RaR����G}��������e\ M�"U��w���śo���^�g�{V�Xo��v���+6�YĐ���F����F�8B��5H<9�]���Z�8y\ k�NM�n�Dw	�v��	>B����u��%� >��_O�����<`[^Y��3�177��!�f(/�b�Ň�?˖-mY�:y����x?��t���'glsZJ�0�ߴ()$�ug��)׉�9� =�O�i*��"r���%k�^�I�I�����C�gZ������|5E�sDg|u���0����Ԕ�J��t�کD{�M�KIڹ�s���?�/xq;��M=��F�M���ʎ��~i\\��b���K��i����b�/_f�e�g� ����X>l�g݈�A�'�\�]SQ*�$%\>�xXUA�T ��Qo�
Xz���ko��(xF����3�[�D����0\j�代sѼ�c=�Q�E\�c�en���Z���c��P�JO�;���g�0���O0g�`��Km%T�7���]:~v6�ݽ�y� '������~�Ɵ~e�/��_ssV?9?�5;��ۗߕ��gߜ�=�O�R��m��m������|4��ѱX�҂)�b��,f;{�k�5�V��.�^��GX'�B�y����=�1>�=4�ٻ;�_
f?����&�Ȣ%\RM��� -͍����{r�,�{�z@��F������~3��HO�ǵs���H���V_#k"k"�d��C�$c�1�}����s��m�mxqjuYB+9���!Ԯ�j���� /�w�&��7����Wu��7K�W��N|���=�|��~�A!���㔿�i_�g���d�1.�i�|��KU�o���K�N�(s.�'�VwWW����yor�n�Ջ+k�F���ӗh��Q%��W,.,EKJ�k�X$c�`Y��SM������7���$[�*Pe|]ͥ�)��\
:�bf�c������Si�@IS@��D!f�l����hn���fD�*�L�J�U��f,�J��¡�Ѹ��K�R�Ux�D%��;P��i���>Gwi3��>O�7�/��3�½��e]�|�� 6Z��5uhZ����XK��	:����z��}���Q��:�f$�sY��;t7���u��imi1�ܻ�����w>~����\��_m������B'��1�<��C�i�Fkc=~�9�?K��ᓈ ��vqT�o���O���Ų�0+@Ǜ�����g���f���u������U�_ƚf���" rS�8P6�Q��gu華J�����X^z�w)1/�W���LZ�}����c�'�V�g3��r3�|��߸%H^�s#��Or���S'9��t��V��&/���#�ˊ����j�k���i�> G@n D���ႥmHx� U���������e[#��<�,���d��$ �r�`k^q�xRW����p���~���>�K���|n:�vx`�x�˘~{hP'�����+��p� x�S��y��Pn�aW��64HDR��'�1ъz��!a
��
@UT�,�Xq���(��fm�?G���f�K�%^o\>x��w�ÏoFskW����_�!i~��q�ܩ8w�/���3���`�����V;��C�N�x&��ू�ո���ϧ?��I���tlf�*Y�h���c����j�H�������S� �X�'����|T�p��>D%�{�<��ɔ�7 B��E@�E\L"�\����x���s>v��C�ГQ%���������|s�����)�>���l����ly��������y;E`OS!�1,;�g�����o|��h�����a���{���-
�����l��^��� l����b�V�T
�g��g����ٖ�K�:�&%0Df�s�E�O��0s�-��}��=,�@�`�8dP�ni=k�ҳ�� ,@ӿ��9V�m���s�Ȗ\CL�M>��t�i��t
_f��眮��z6 9��u����� .T�<�S��-Pu���n�V��w���"��M�h���(U(\�v�?L�Cb�1��4�[��ˉ��݌���<���C����U�
�� ўv !�WU"	�I����0)����$����+-�'��2033�#�uPheU�#r�{������Ac���p�,A-*�	������hϠu�7�RJ{WLHSE|�����W�S^i�'�ۇ~#ʭ�w�ɿ�"m���b�jih��m��^Z����q���n����͚pJG�B�0m��Ȅ��2`콮�hY%�}���5e�i���\?L:x��I���S�)T�x�^R'����pV�y��^�;��KfnR≙2C��WIT'�!-[��הzà�;���3�w4�����#�s��~�plG�����������J�~sݳͿ̨���������տ���ar�d]m]�<uJ�|�ۘ�m2����	���N�����R�Ed��  *�D���Z�xC��i�|���`��9Z�!�;�#.���AR���)jIoV�x�(3�*=AyӶNǮC{I�`�(�?�crE$-zN�-a��
pg0sk����vw-ɂ��(Cr��e�ֺI
y�h1���zW^Z�����O;��Xz`S���ᖬ������T�UD�y�-�=�_�4���C���Q��R�a��&_�b0ϩ��r���� }�'�Z>�|�� ����a�m���g�&��wR>+����D�,��*�ޠ������J0�N�c:N}K-إc�>���Rv�OO�v��h�]��Z���/��{Iْ�R �U+�?y�;._<�.�qOSJa��}eRS9�i�����pxI����=����P�4���$I�X�ޒ��|��P57�:Z�Z('�s ���F��!�x+Bf�Q`~���D"�Ì�OO/r���)l��Y/E�w2XH<.�O8���~���f����p}I�������N6�F*�Wo*V"��n���g�,@�>�4�@���7��X:���p<���55�b�Vko��ǥ1=�c+'�&�'̪��c�/�'�Lw��m%`ɩs�E���8�ǭ	ERF[&�4�!4<��]9�y9聁?Gz��7�(b��Lua%���"C���E۠_�],:O��}h�;�բ�'A�c�K!�R��򙦕�|��|�Vx/Qu�5����F9x���V��#��#����4k��]SJ,���Ji�\9O\=�*B�h`��2P�,*���r����]X�����v%2���ѿzK,�;�:�K��\�5�dO�J�>����=�-�݂5��P�ۂr�'4D�8{d�1��S�۲�5���Wɽ�ޜ'e�����YRE��:��^�yt<�1q TE���",��Ջq��9�6�Uy���i5OR�{��H/�$	�H6��LP��U@�'� 4~ӭz������r�_1������ �Yf�qy��X뗳!�-��?L4�N=C�ff�\�Fac��k:)1JJlyU���eP�E��3�M��4k�������|����+�WoT�k�H9�X�����N���y�ئ��	���>2�����c	�q5T�y� Ʋ�{����/G��;���UѺ4L��ݼ��z �p�9�D��L`x5w] ���t]�z�1!�Iϊ&, Zݏ8PN`�[���s�"yp� ]<�>� ��x�R�PV[E��傶�I����y�S�������1���퉠a�aB=�� �e�}�~S+l�9?���d��}W�
��I�N��3Z<���`�_
Y�d�`�����tP��M�*���cM�ş��wc��p?�����p��?�2�PgF1Kx�Y�|
E��,ؓ�����sq���h�WW3{[R��-��?�ăvq	�/l<���lo�R{s��6n1ޜo�Sy>�8��
�c'J��d�l.De�^�t�K��Ǯ����{��^��
%��A��).	/3:�K��Yr3��Ov���<���|�p��,%-�Bұ�wHhu ��G{aV/�T���e%"H�./fع����'��J�thdݝ�j �	흦F��ZR�|���|��S��F�ܖ�.��(Oj�:AL���t���?n���-��p#�l�����w����~��Ϟ[j��O�y��O��58�aا�5�.�A��Aaj"f A8\��zOFY�$��\YF��ŊL9��l�L�!#Q����5{�}(���Ϭm�L2�q��� (�p�����d	�-_��pѵ�,I��M�<�s  M��u���kkieG���ZD-1Cس��V�'4f�w�e"�'�1ȃs��{m\|d0W[� ��c�%�мq��:!j/�S���n�.A³D9���ޛZZ����_-khj���ƨe	j�Z6��vBu�4�ONDsr��όUk����v2S^��}��w%$v�o�U�Z]��!Se�U=�،pa!���e!p��m��64�
�/LNM��GP�`P�H�����=���!Я��+�I8�=�P���M����yac@�[�?�S٦/Z|��<�����tK��W��3�lBH����×ܽs�c*�v\8��>u5�^9�
I���t����8��>*��`�ԠTT�ԩ�zV�������0�cߦ��U�Dϫ�94���ٯ�)O���ﰴG ����_H���# �@ �mE�O��;�<B��x6�@���[3@��"\*L�P�f#����&v�"��o߽�z�T��d�̿��9�7yz�-�_�ОD0jO���~�vVB��V��Rn��m�?�ْ&�S�������O]�}�y��3�Dd0�&��R+ؒ%��}4��j\S.�oݲ_��*��af�Tݱ_ݚW�ؾ��Z-�:��I6s&�D�HDD&0���g?�Cv�̝�6������k}��k�㽟'x^�z�(C��4�^�ɡ?�����������*Vٺ;�U:8����СC��`i���������@�mP��Y�`i^�0��4L,+Mi���r��������&e�M�@��f������(Q o7m�8��Z��m����$k`8��K�S�<�w)��+�kJ @B�|�H_�߰��A��ͭ%_J��:^�6�zJO���:玹9*_�j�2�����E�t�މyfZpaV�Q�\Yh�,�Ģgd=ǚ9T����m�+ w�n[�[B�2��w4c�VYȨ:q�@��M�^�2�X�n}z��˲�1�M ���5Eg6��ѕ�o���]5���F"���a��T[�C��+�+fj�
���}e�1X��3
V��[��2T��O�j�x��8&\�1
u��敊�n\�0�v�aA�}�X��6۷��X�tX����
 � �r�h��!h���00M�,���͏��+H��!x�����4��ա�o@465 �؏�2�BUT2�$��{$Y�ߠս,�eKw�kشyS��XR'O�H
�b�,�Ֆ�Nm��@3`�pB��m��b� �����q?�/�H]�{ǱG�2�[b�&W(����k|�?��G+�y��ſi����ʗ����;z�EǄ46��E�N��?W��oS�l�P���e�Ga�z��9���1 `������_��U��"6@뛧\6���e��EִMm��B�<\t=Ѧ|e�+c�"��͢�jf{�y���q���������~Kا�@}"��.�[��!ǀu�}�3@i��)��SP��A�[��Z���n����Fs�Qp�[���(�i�b 2gΊ6k�Ԛ�KCo��{�E�>�8�f�X��Ē��q�O/_�_:?�LۮZ��v�=2���b�_ �ҥ���^��3��H�/^�,������p�i�g�3j�ea�3l�����w�c�-��7k&� uV�`��An���Jv�"�>K])�©���]�~��"2`NA��"�*����|��bt����)���j!���
7���{���a��5�������m����$S�݉��7�F�7Y��C���u�*��ݫW��&3�lv��zn����m�=�D�g�i!Νwn����AlK`��	�����U(]�!�o�O�7����M�I���+���k�S�N�JBZc}���>���M{�Y�J�O<�b���O����-LI�3�����������|k״���3i��J�щ�]۔��%���h�۠�7t��@�^&�j���my�k']@4�	�+%�h���Z7Ǿ�Z '�m�*�Kʛ�#�3 ��!��c�ܥ��e#3G�(^�3y�hU�p~�_��X�OҪ�#� ��Q�z�ʿ}�Jݽ'({���$V�U�M��^Jk�˭�vh��ڡ�r�6Ճ)�������ǘ,Z�ϛ7j�5����B�y��U]�C}��:�~���6L�;p�KP�5�oʩ�4֬^3<����-x	�i�MD�1J_[z7��Ϫc���E�L9*K��������y���?	cӆ�˗�R�k׮���7���.B���o���5ɹ��*�2�c8A��y�l��LIi�%�ʿ~�� 	�4w�Zz�)P���s�F�S7��j������[$�q��૜�u$M����4�:�8�Xf��K�@Twt�*�T�w�r]�R`����7�G̹t�֞S��F=���d����3U�^��[ʟy��>�F���?+L���>y���&��R �ҮS��i<րE���b5)U�A�{ڽ[��k.�B����n�p�Y� �Y�,�kåX���B���@�ܽ��1��OS8��KVr�_�����V^�$���Q@1��I�g� (K�l˰S��?�W.`H导]&Ѵ�ɵ�Qټӟ�ϋ�����^-.C���5��ƢЮ�yp%`�2n
[�,��=62��6�7Zv%��U��X<�#��l&[0r�Ѯ�����Nya��`�C>X�
l����k���bU�p(�c��7;O�g�0�*��5=i�~�z���b�\�ڋ�I�ݛ��j4�m���h1਀��BB
�z�B#"h+���D���њ�L�Y!l��8�_���U�*1f]`3�J�]���>2D�^�˯W��Z���M�ڹ����ʕ�k��ն�Z��n�k�e�`b��7U�)�|[T�������ޫ�&��ڻ�z���N���/'�
�b��9�8d=�NS��q��'��{}~L(Z��,���H��D�V]lVu�3�K�г��ϕ� j���̮��>����x�]��4��4F�G���f u�`��w�;X�C�_�IS,ei�9&�*C�r���$���g���O��`����3v�c����!?u�j�LͯoJ��� _�����
��#�Zxm��E3ej_�Yz�Ґo�I9kr$��^�N�bm�lK���M�5����Q�&�ޅ,zmZ��������Ǫ}��\W~�?��aÆ���;�V�ʊ5���*{���j�nimc#�=�H-�?�^Oz`UwkOF�(H�������?)�_��44�+,&�B�&b����a���q�	��0bU�o�ʳ�1�1��Ϋm!�S}���J�s|����h�`���ۃd�H,�wY��L�[W)��/�[���k쪛�US�RUs�-���߿ic�r���LX���5�a�7�?�P��t@��)��9��^����􆝌�1�4����=L�^������,=~����,Խ�?��ĕ�-���۵f�7z5�v��FW�S�R�(���C�����]��5@�j���ּ�؀e�����%cD�߻�dV����R�[Zz�N��+���_����(�:������,��7��ך�/F��]�|~fL� ʒ�,�Q�N�h�m�@1����r5E֬|�t���ӧ}��m�^��rT�u*D���JD^,ߞNk�mCWr��;���{��r9E�K��w�|6�\�~i7�Q�{%��E3�r�Y�&���m]z����7�M��.HZD��Ѳz%�/u����=ݣ�k�RaRb��Fc�.G�>:|�h����z�֚�sϕ��
6%~�9�O���_<�p���'��O�iX�o��^�Ī �;y�1|+�B"���L��p�B�=��)M�[I��	#�H�8�(�\�J��B���[����I �����nI ���<y����+K߯���nO���Q�5t�SS�lpE�P(���ۉ�OV���ϻ~c��ޣ��bF��-K��O�&B#D	�D�U@���3�?+ �ψ���؟����gkO�~vh S/N���$[;���>³v�Ż��t�HỲ8�*�e�����Ey���n�6G�4�[~��>xO�$5+%��J(AMZ�W�[ 3�He#M�'v�%�q3���3=x�@9� ��kr6	��riLI���3�����  .y�N��Z����������h�k�=�y���`��Vz��V��^��#M���,��ʒO��O�h_yً	��*
�J��׶c0����^��Mo����b��۰��<��#��-�Ӷ�17���e]�6�)��0~t�K��R�P�ı~��W������/�{���w�N��`QMi8v�Ќ����=y�ǉ�4������J�:�*T�P,!L���~\k�@�Y�]C���m�%�g��VHsd���wx�����{n8���1�4�qK����و+4FDӖ��x��x����p{C� u/�fox��SN�TtM唽r����i��ʪ+PNs�\2[ȪR��޻��v��|���
���Z�/�J4�#�.��0c�$��˳�@�]o��7>ӏ?g��ϊB1tb��ri<1�[�J��>S~�34n�������+V�����*$�x�����pU6�Qi'M� ��J	q�_��j�Dִ���f�\����V#� mT+X�X,�(�IK����e�ү�O�%�JY	���<�O��o"�x��%��~JL:%��0�_����$69�rM�0��s�ӿ?�^���9W���+����N�x<������o��G��z�^�P��@�](G/7\��ߌ�����L�h�k�M�qǺ��(����*�V�6��Y�?��N��*cbaDx���W�]�d������^�����z�������7=$�'u�;��Z�I+:oA��8�b���?��CY�F��B�W㌢�
׀�ISɺ�{��W"��8r�pY]�Rt���Q_2���Ǳ����YD�Xa�}���~��p8����9w��/����,�u+�J�d/g�������^+w��Xj )��/�����ʌ��rջ�~�6a�$j;�4�Շ���7��~x��� �
�u�8'�5�֑�J^� t�O�X�^�����C]�l~�2~�����0�Q|ш2qM�h��Q���$?�a��ʊ�����v��KG-�l�N�K�-���jj�F綘�ˆ����:  h߿�����Ƶ'b�j H����V{j��^�Q���}N�ud�d/ _��BP��'O�'-�r	h��� �(gb*�7���Qzʋ�EiT=����v=�:�z(���t�=�ީ��k�����������[��_���K����L/�{~�_�s 2$�c��2�v�/7Z9���ŋ���c�fp� u4�N����wo�5��2&���Y�7��v��#-�)+%eA���ѫ�Od/�)���O/>>~��ξ+r����X�����u�)�ֆ"������L�-�t�������x��I˲W��Wu�=�S8�޿��ꫯ/<����~8��������{��^����l��@�Qi�Y�|�bO��{��OO���klA94XU�����A��Em0Z!�c�K�6-ܬ��H,F���<�a���~���b�Z�gru��hSeI�p ����Y_S�l�P������.�;e᧼zH��BI��8�����կՄ�;�2�u����?O�$���zxij��v�����Q�N��t;�泚��Λw��/��H,���ڂ�f	 �v�����n ϰ�k�����w,�z � |y��<����D���_�s4p^S.�E)W[��!�����x��),��r+�n`��+��q�-�=5Vo��Q��5�!My�M)��O�0�3�[r��CWZ��eTPO���Q(�pϕWY˻����;��w���g�����HDsF�ɓ'kmj��t���V���]�7�˻��i�C��{�����x�a箻�^��J��c��4�CzU���s������J�=�k��Q>.�E�n�K��k֮��K�A9؜Т2= ��w�J��
+�eКK��!��X'=�t�������� ���ݫ��VP�Z�o��X��������x�������eI�F�eв�9� �U�M�Y�o��[אַ���4��tw�>��Puo4l�OV[��j����b�0!�D���T��X	k�b��P���i��$_�bY��Z7��>2嚽E�U�k֬�&-�DI���2���&��U���� w���g�>9*,*��S�Z��6�[��y�D;'T�?+x�+�������ڔ�v��c:��ڍ04�w��`�����w��)}���;! ��y��W���|D�7���CPY}������,̲�"<�4p�r��e��*?H�����;_��1��{f�h[
ɬ1S�mK@)i_��+Mz&�M �ޣX�H���w_k ���W�"e2&��Q�溲3�o�gi@��Q��W'w�WGۤ�`)�i��*W7vZ���"���/]`����`}s����R(�^�GS�-������E�`��L��H{��4�?̨i�^jmPӲS�3���v-0Q�e��hɝ�٩�陾p��r��'�x�>�nϭٳa7ϧe����^*��R~Gm�;6|?��o|c�ַ�U_l����W��^�p���å��� ו:-�|��h�OSI�����;j��a�}��o��F�ׇ��z+=�R�[e�+�,<p5y(7b�{@�(t��|�-К���=��T�ٲ�֮Y[�����{v�����m���I��й�0�=s��b���1lj�~Æ���-[�-��#,�O r�5{��?�������G.�c���������(*So'U�&�����(�|�J���\N�`�Ux�~+W�RNB�b�>�F�=��%K�Bc��A�}��JS�?a)�<:[���H�(�E&��Y;"P��@��v����&J�ݔ�������\��﹖�~��쎣�ˣ �)D�Y8����+?���f�G��ʥ�	):�������0���w���.x�D;�j'��P8ڙ����g��k`0 brA1)���C�]H�X~�O��hH���E��]�;Z������+"c���K�[�,dZ:��Qt��Q-{�,-��x����C�]�s�OGͣ<|��e���2���~�f���mQh�i�0�<���g���H:�S�01äﰦm��]-����)��WђU�%�Vϡ�O���J;���m�޽�f���W������k��KW9�pHY�,?������o�#_z� ����������H��� 7\c�S�f2xF�0 =�����6%�R���?�P~�hl�AP� ]ʩ�������~���-�s���s�|��߭}����/�����O۷o/%nܸ�a����{�鑇b�#�� ;�WQ���'sr1�};K+�o��d�f|Ϟ�4�V��ua!�w	�t�M!k<��
���I�V��h��4�jD�с@~���`����&|Z���{����ԓfY��ħ���&���z&�1E	)o�V�E����V:6��E�4Я�ۿV���0�����1���k�)�~F�4��G�Gp�s�����+�~�p��b~5�ڟ�/�����EPЖ0�Yi��ќ�.�Z�>�pm� 4�����W�������Z��1y���w�/ >J�[�)�rK����Ʃ.z����/hsV��� 0~ʆe����<%��T�(4��dC�kI��"Sm+�(� >�f��x�s����+�i��ɹ���I��S�QP�z6���,�7�J��mS_A�}-�;ځl�����*2Y_1���z`�.����LQ%O�8T�η�E�-[��v�,ctָ_������D��;w�:��ª�{�(f`h�;��[�s�y��Ý[��vSޓ#Qҁiڷ<�M�0@�����Z���93�L2 '��o���[�����n�a"��?����:����DUH�<X �n���ޱD�ǲX����tM�( Z�uc-���nǲ5�h��fYD�/f6ƵX�,n�A� �̀Q x4[�#ebMx)fq�7n�R��mSK1_��M���j���jlQZ�А�$1�@��?g #A�ڂc]n�s�����;!$��6��sޢjL��]���&T��z��ｊ����E���=��c�R��Hc�VO������Cd�";e���8}h�|(�E�5m��J�Y��U/ ��*��}��W��[(( `�2�/���G�w�J� ���qFR���cz5�LXz�Sj�Gd�ה��e7ĉ���7����6�$���LSl�c��;�����EVfY�9c,��+E�G!ځ ��4�S(����x�&��
uo|.i������v��g�5D���C�]��\�=V3���Ν=W�*+��77��<Kf�w��L��C�H� b�g��x#(k��g~�o���[���ï�گ��+�2�����������{��������R�o��fM�J�g�0����<������/������7w֊��(��l�B�ھ���|IѲ��M!�0����[�9$4zL�i��!>�����02�	#�@j#���7��놿�����a���iIۗ4��L��{���K{J�?����}��7�sϽö��tm		����bSJ�"!�|���h�c:�������t����#ñ�����m�D��
P��(���?���'��oQm�,c�-��*?AM������B�|~W��LP�$[��K��P��,?=������d�?;���H����ϔ�?�!��Ҁ���p�%˖V������K�������Uz>��+��3�F�7n,a�̾�����[�:��|�����	�C=��4˧͒;g����<�:�!�-�b�7�l�?^�<#GnF���yb�g�!�L��UX(t�,�6`܁��Y�)0��u�۷ow@"��������Uco�)�DC�U'���ߺ�R���A=��*6������{s?c��}�Z�9���ymV��R��js���:jw�Ѓ{ ���(A�O�{����(>�����8/�h�i)Z�܏):J��;[9<p0�M+����ޗ��r����h�\l�ß��|������b�3t�q%��7�x}��?��z�W^)~G=6��)�Gytx�k���tʥ-�6�q�9����в�	M��6!,��B���j��o���h4:!;�{|�a��s��_�U�|h�Gy�*�b(|?�1������������e�];w�?����wӍ1h�Q��n�
�x%T�s-H�8���:���,�F�z6���]0�ޘ��F�K��9!e�JF��y�F��L�M�:Ϗ�Q���Si�\5��n3 P�. �wZPZ�>�<'J�sD�~lr�z8?W�~��ky�$�o�����7ӡ���3*:�7���HԞ��%��8�ڣ�U��GX=+�3,��\���}�x}�� ��ǐ���J.�I�E_~�+� O��,�k֮��;~{¯ݽ�\�s���b�Nrlg�m��;�
�K�m_0� Z/��lK��Q�h%:�n�}�S�)�y${�'���:dG-�~y	rT���J����+�4E׀1�EVᅴ����m7(k��升j�&��#K��ћ�>Oݙގ�&7�O�D��R�����=5#L����@#���y��2^�|"����:|�y�RF#�y���\��
���ſ�˿���o�X�V����~���_�Q,�DIm����
�b��2���0atzx3B���$��3A:Q0K�M�W�.i�KW��k�CI�� �K/�8<��5ha�Z�&~��Ǉ_��_J�u}i���]��?�����zF�?��C�c�>6<�������kpC����J�H>��N}��W��ckQ��6]��V�,&��1�NQT�  o���Y�� ���x�I���ʀ�����B�n�(�sM�|���d� �W ����� i�Z3�?t�6���*�v�_��s���&Қri"ߟ��hQ%�^�O��6�{����� �ϩU�r�:�^T���$f��Bl��5*O�_�J��P3l�C�|��J�0���E��:�v�em|� B�@�a���Ue���R�H@�(,�io�SJ 4���:�.b�yV�W��k�']��]�����
s���~wO]�8�' �s���}����J/K�!_ ��P'uS�ܬ�_�zT>�i@ی%���3�tsT�m��[8�KQ5�l�G}�@��E�t:6�܌<]N�*K��m���$���M���<ԃ�ږݶ�Ҩ� )�-	b�3��l��\~��` ��=���ʯ}���e�`p�K_�R�5�{���B!16�ʢ�/�x~��fu�5���50��/~��=�V
��%/��#�gCT̅(����aa���kv~��%� ~o �ڵ�
�裏��Ҡ,��G�KZ(���OD9�w��Î�wk�`MiqJA�c��ԇ+R�>����XHF��۩iy���Ƭ�����x�NH��ed�< |!C}�5�g�Y�H�M�`FVd�1���&���f)��&]�f�L0{2-+mLmS�Q�[YL��u2�IQ%���Dۏ�������G�(!�&��g�+��)�6�I������\=�����\=K�.@��{�Ύ �riX8��/�N���=c���ބ��k�ٴ��GG��WTzF��Y �m>��L:����O���
����*/ �(��6 �M��ˣ����<S	<�~�;q�S.���H<R�y�ox�Hj|jC�f�;�����o�oeFȋ��ڱ?���]�]2�w���J�G�Uu��9Q��8�LR��w^k=�\��9�zM끪t�|Ro���]�r�Жr!o�M"o\�,Ϯ�QS�h�]:֠�u�a[���3��λ5�����^���۷�x������XF/�Sv�tЀ���s��R��e ��U����B�T2���lzvH���[j�@{��5���N5�F֕6����XG��wP�`d�wz0ZJ�XP���h#�c�_����#w���ڲ(XHY�*W���U�6h�K���|���QBDڰ~}���2�R��PL�k�����j����X��_��ao�>^J�%�A@�>:HR��r���l��+w��6K�)%�	�O���Vy��2�X���yZ;��ڮ����(��K�S�U��i��=1��ԐK�w~��}er>�\b�Cۅ&��w�g�r����mX_5U3�@�.���:wK��c-��k��n~s�,��- �^Mԓ�ɯ|*הE��s�W����' Q�I��c�nڼ9����E���e1�{���2��\���9^���/�EI�7��#=�_�T�P�^�j��X=�ʷd�!�8*��"�Ǘd�=e��{����{�d�u �����<�/Y���a��Დ���]y�d��Lek�Pڎ�\9 ��R�	ڣ�����
U��5�޲yS,�u�zd�������{�ý�oxȫq���Oe4s��c�p6�t�@��/<9<�ԓ����S�f���l�Z�\�6�L�\�<�Iz�[��և����LV6�=-����>�[�^��?�q��s�	3�%��#���6��`D�%m>�-�ix�*M�a)���^��E��f��#�p��-�j]%�;&�+�(r���%�Xz hb�z>�R�S3׺��q�M�b�4Eq�ʵ����a���g�Q�X ׮�y��)���+'�X{�l�� ��.iy�¢	P���E�r:�/�M��t#D��B�Wʑ��54���)O���b���ޖ	�>��\:uZ?��.^����C�:��Z�W[��q�&3L}s�F�1�
�]ew��vR�n9tJ���7,cGg�Lq5�����f��ݥ5��k�\�{�\`*�7.C�&���)mB�S(�}X��m.�qo����'�#�Pϥ�<���LM{f�����Z�_|�4;����u�}J����ڢ�2���$��!J�m�%��֤QO�����%D���ԋ��PBJ����jڶ:pa��zp�h3`���N�#�K�xw��j_�.W�:{��-��FVE��-�OY��1�����Z/;4e�C�/���
[Dz׎���_��� ���~��;��	��,�|����󇕫V��wY�z6z{��������M�7Ӈ��F�}ʭ�t`��?����#1xl�cl��R��ʽ�:��0����2����Q�ot���8N����� |��}�;�����/����R4�˯�R>������;����þ��
�Yb|��V�.-&����w����_�~��t�^+׍Uo�({�2k�B�r3�7RC�K�г�>[
����[�������ؿؿo_E��E8o^[����)B��Rj��b�rτ����!�,���X ,4m�o箝Ý۶�?��t�i��e%�]��0c941|O�tˍC�)�� �h�l9�wE��6��N�Qa
�*��4슀e�zi���@���P	�O �YLX�M(���}+��鴣���U'eF'�������n���]}�.�I���}�!E�i�st޲uK�����,��]V�Z�R�V�O"�+ϊ�(Nʁ`b��>�K��m�Q/J��,�6��f���`� )�.]����-�W�w�xA/Q/��z�F�F�rI��b�V�$�n�߶'*�
���{�n��^���S߭6@�\�V����k����-E�;�(N42���Z`�> �|�fB�7��3}p�&2�y4)=e����F�/��E��������=�X�S�)=�R�pl��#��{��R >�(\������H�eX&M��\̹r���Ѭ.�P�?��b����z��>0�N��3�_F^巾�횾IM1gd2�_y������χ?��?~�����Z͞To�f)t�Ʌ�ed�=���}�����tfB��ҋm�9`��Y�vMUD�����nc!n���{7�?UV�B��z{��3�����^K�?:�QT9�|�����y��1��ۦ�5�7��FЁ��{x�|�ᕗ_��pQW��(��s���L"�&@p�s����+�8�A��G!|s_�HH�k��d�6^�|i�FZ�����<�f_��} \�j(�#�#� ��e@��Y5�2�j����{�3�[�c)TBF'Є��T��G�;����5U-��`�2�&��7�FW���?b1�=c���2�9�9�T1�OUiR_7������X�� �n�w-ڑ�p�z�xI���̅�?��\��jSM�C/ϳ �E��̀�fI��˯���ݷ��ecq���b��wY��>���ڰx 啎����Y�������� ���y��#D�F��_�Z�����S΅�K��ЏE�
S��s�~��S�7ۿd��RO��3�~�!�z7m!e�����
P�p�|�g�20(R< ��^1�����_�P�Cz����g�DϜ�6������n�k�ed�{
^%�í�7�Ӣ�6�`�sX��b���S��땁�Ȼ�F]o�6ES�OԀ����jҶ
�S0����¬(  ��IDAThya����?��?)��b�e��l�#�ٵ{�p*xb�?��?�z���7�f7
�:�
�y���+"7��b)����C5�d �6S����_�����?��c5��w���U��׬��Nf@ڨ;ͥ�uO��y1�ҥ6V`PW;v�H����/�����J�p\;�{�? .@ѿ�V�4�A]����U^��>�C@��j�{ұ؆2*����0y �h��1BL�x��<� �Y%fpؓ����ra�%���ɲ�i�,��|Y�7c%��=�15��:h`�Y	&ꪊ���ӻ5^P�i���X���-�ՠ>���d
��0����Kdz(�����y��CB���V<��U��xA8�jV`[��}�C�E_uU�Js��n�Y��U;?�qҽ�v�|��<V�|�?K�)��hZ��E#i���$t!�5� ®�F�h3V�$�K���n�l��5esT��T�u��i �g��|,:#��Z�Y�]�'3%L�cjZ9�<&4��1NZ�zlT"�A�k�&�3�Ĩax�S��s����vt��s٧�1&��G��LG��A[�e=-�!�Vr��f�.签�����:����"6m�P����d�&�xjo
��9i��x@��4�?��?��
�������^*�E��p��Q�x�%�gX��r���董G��|�;�%1���5��d��Ǐc��.D�RO�tc��&��
>���`��Y�\�U�������t����Qb����;���������X���i�F��lӔ�{g
���L���-��#ټMe�,t���J��3�~m�28Z��<��9�{۴is͵e5b,�e��3)��)��5l�6U��v��;C9b.'��>���46��j���D�@�}e��t0�|�����%�<K5 �=�1�eΚ	����>0+�Mޓ�PP0��b1s�Q._r� t LWS�����%���[9�է���ڬ�UՅM[�k�d��0�ϛۖ�X��Y�R��M�4��-N��er��Zh�Mf�H���f�LPo�DF �V�&�3��i�Q��k�pW���63E{S �D��{�s��^NJ�t�Y��	�|8�b��=���ծ��J�x!h��.�{(��?��M��c��3���Kg2�
�J"����b���MIU�-=<��V{�s��ц~�E?S�����˻�7�t�#<�g:�#�m��v��%ɇ�0s��O��NoB�ӔNS�����s�jR��N�3c|n�n�7�?��ű�ɕt(6�ki4���kO�}��7��}�/����=��S��W�n�/7�^�fX��:cپg�1#��W_lCN�fj��o�YE���w~��m��mfKyޓ�b8�9�e�ᡏ�8�O<1<���������oW8��m��?\�Fʲ�B�p]"�L��`--g��f�����>��SU���`A#ύ�_�HW{Ir�y�z=�{ﻯ�����_W#?��C�����YBQ$"E�h��h����k��%}ۅ�85(�{�p%���6�@�86��{A^`�tɸ�΄�ug1��{�@!�j�@���.�%����go�K�pu����t�;0�O@�C���0L��+��>,��c�=OM�R�0��ʱ�08%j:!���0�/�e��A4 E�Z�?oN��R��߾����X�zy�{܀���c�}�.-Dٰ~ذ!�B�����r޽�L��$H!x� ;��	�p8{~�5���?}zS�k֮N��GXU�֔R끘�ߦPZ����z]M��U�厈�+�bڏ�R���#� 0�U2Q
$��y3Xl{����vĿd�MS�o�\�=N��%}���J���V�ڵ	u��W��]a�}�) &N>�z�(/%���^�[�-��-=3�6�ٓC�i&+�ЀK͌)����vAC������{��O�3�Гb�<,�ކ�����q���#���ߺ_�2M��� /p��0l��3��&��lP��t�o�*g����������v՝K����b�=p��%�\:�#�|��2x8�0��]��k���- ����?w��r}�:ʂ����X=�@p�G��-��� �l�f�&a����7���o)���j  u3�0B��+/�
4~~�g�VMI2�y8>�W_{��\M��D	wY&	J�[���F� �#�:��(�jZՂ���0Ƴ�� A�+������j@��)z�o�O;yM2�f��	#��qB�tY!z8�8U �B��������%��Y���������K��zbh���?����Սe����_E����Xs��+���W� �(pU�o�2�������=��#Ó�逸�0|��O�?�h�+o_�.�@�t�3%l���j�_��/_I�_���_|�����������6�����沮6o����<�z��J�}��8M}#��=nY�h�E�6�j�i�7چjf�hO���hm ���k���(�a���i�^�r�W�@��g
�ۆ�ł���+#�_ڵ��叒j~�V6|��u�xn���>`������F�����6zLF�1��;NM�賿=)2�G�ђR$W˖-���. 7xːQ��/�k�2���_��ᢌ��Qt�}A>"��6���켕M�W��G�t��nul�(3�z�u��)m���M(��؆��i�娇���j�rikg�ڿ��Kep0x��r��Xw�&���k��VJ�l����;
�Z~��ɬp�'��-~��1�ƒ2[������������K/�4|�[����oWׄE`�˗���_�@8����/��߷�f����y��T���ќ��:��?�o5�G/��V��K:,�w�}�� ׏.f`=X��x46��zA��6�`�"D	bMc�t�ӷ�d���Ѱ��Yh���Ф�~+SY�W�~Ř��N���]�=�tk�y��m�u���ý���l�B]�2�o�zt�X�f�@],�V�K�,���w�=ã�<<N�k����%O��L�Qh+m�z+�n�/��s�ܳ�|��sŊe��z��\���Qp����!�m�vg�my;�߬*��Z���Щ}-�,�x�z(�?�h-O_���V�
���0�t(]]��mŤ!����l�;��з�&��Ɏ��* !H�����$�<�C��#�`�+��P0e�VO�Xvh@�p�@&�[0���S;A�)<�����Ǐ�J��Ty+�D�	t7�Z~�lϻ���������Of�ҙz^y���O���z���ٔn{�]c��]��S������i�g���^=+���I�p�:JX��gFM[�o1e�(S�4�/#���k���Ӗ�Ps�o�rP���˥�mR��������U�w[c9Q<�w�o��}x�6j+�<��yX�^|a�"�� ��a�ј���P�q�p֌D�0����� �����>׸~���_*˞Rѓ0C��*�O��?%���
#��PjT]�X��ɣG۲d�R�0Yj*aN��_z�V�a
�FhcY�!���6C�@*�~���霺q}�
����FR1����Ƭ���_�ձ�� ������1�y������Y<�g�4�l�z䅱�a�����5�V����I#PP�BG��llQm
�ڵ�"sfU����l�ҏ�s��^�@R\��\=�"�=�H�-��Ag�U��@i��I�s�覚6Ǌ�7������Ċ�j��;��5���'�,��+023�ݹ�ʽ1
�����4�� �A(����"Di��Ҕ��{u���p.��4�w����]�HM�d�Q�,��6���)�uw�-�
@`���ztxʹ���I9�CYXTzƃ�ˢ=�S�X�xѦ��#�b�^��\��,hJE���A�π��n;͏��Rcp?�N�����&���PO(��G�g����)��Ɣc{�}S@l	%[9W&m����-���7>k`�f�Q�FW3{O���U.mƅ���� ��C���sư��oM�~��[�n5
O�i�G�K�)z�XVw���ż_=�J �K�e��:�ҋ׻��\�f�.*�LkG��2�� �:�n�u���?d�/5]6ugTuZ�W�e�� �I$�/��`��wS-n��6Q�IP�Yɘ�������[�W����t_X~��Br�S��_���o ����0%�ц\��;�;��/}e�'��B2Њ	 H������o��o���|��e���<�b���ಡ��R��a�j���r(�m@�a1�P��н<�許�oְ�.Z<�[�~X�v]pq�o����6C��\T���hi*��Rʏ�e5��Ā�<	���xɗ�0#d����0y��K���잦�
 �+��!n���nk�.?�ȯ	���o[�H8��
�����0$x���<���Ǖ�д������d�N0=��LM�MyL� �����
@�')K�Twc�&�� -�����`����xFZD�}�/ �s���k�)��ړ�g5�
�k7�I�M<Z��oʮ���N�1��t������~V xi���c�?Vh�j�v^O����'��=(;�[̈́��3�+wG�ݍ�6^�g�~�<$�1ߪ�R��Gm�6EC�{@/�G�kS��,r��#�r�T��ɖ~�%=����P|�Q6�l�X`��=�1��5��X`��i~=��P���Y
�L@��ofK��o�Fm��y��_�������<����{�-E��[6��w�����ra0��8�ͫ���S,��P*��WA��UX3gʲ�wﾧ�ʣf6`˟�=���WT�m���o�H�mظ�^��w޽sص{w-~�7��c���!}�k��\��H���)��|z�K��G1h��T�'�4$�D\�\�f�%�9{fq��+�k�__�����n�U�'��p������K�-��V�X�z<����sZ@���n�M��q���s^�n[��ȗdΔ�{(=(V{m+�� �h���l�Ɋ ���ĺ�{�cT���t����vw��6'o�p������+�}�X:ɸxA�ô�{��U��[�����])����}����E����2��?���5�
}\�H|�Y����;:��3�\E ��zJ�X
��nw�H�c�Ym>�3���G?*�7������v�'@I������%i���n<�AOD����].�� _-���Ċ�0�0���ej��ϿB�1t���F#g�	���=��0�'�,�O9�����۳-�Z�깊�kFR�'E�} ?Z�7:1la��:�+e��0�A��?��j�S��P����?�C���4�ej��QҰ�����۔\3��B�*F��;�5�����=�z�.�<���7�C�2RJQ6�.�Ĳv�IoC�/�~��`ܷ��A�W�g���0�fC�&㆒���b����w�w�/r'��n_4�ȫ��g�[D��-���v�_�U�'���f�P�5˜?�@�L�ȇ��iq����i[Pg��$w�m�
�-���|5��4b�R�[O>���o���U���6K��L��Z΃�+��sR@Ǉ��ÿ��ÿ���z���_�/ß�ɟ�b��ǎVW�"��E�b����3�5A�1WCc��S&�@ε�L|�m� GϥR=���)���r��Ϟ= �8�>&����O:7 ���q�n. ��Zz遤L��~S�@�f����̾\����,��I����\G���S������?+����ך�k�5p s,%�w1>��^��BlS?(S�*d��8܀��Z�@P�nx��k�?ɘ�*����f�ȓ�M9SN]9w =$��ژ��<q@L�IOY�dMF@O�Ŧr��}�=YP�V���~�U��*[zj�,�KJ�D��Ֆ�,G��N�Ɨ�Y����FK8�չ\�M�}���t����O�EϹ_4���zOCh�J��ގ���(n��3�%���u�pc0P�@��f�1�����ҡ���i��^�K���'fT�9
����&���ꄗ&,�\�R�&綖���e8�򉱓��3z��9�ֵ[51Ř z�E�p~�+_��詨)��!�����S�瘒i�G7x�q�f�J�¹�M{%{� ���^M��E�
��J.�������/������?����o��FAk���z��F��0�@4�g�g*�b�:�����E�43Ķ� b���'m���
[��0���s���N@��p=�47�x��1�h� �oN�ռ,^-,��t1}YV;�̄)H`��_Lo"����[� �}����L+�[�`��Kc�LLS�L#bhS�	��^2��V�u���L>���%+3�9z��feQ^>L������8�a�WLB Y���Q��z���Xm'J�a�8�t,֋�uB$X�d��o�Uc8Ă��);hb0�o�R6 �@��{�N�亮d���q�J�=p�}a��^*WL�5��o��0��:ڳ�}
�\�;>S�X��}��l*aV%S~�eS?<����Q�<ʠ��C�ʈF򑮝d�9�  P�e�,���j���/����]�V���gBؤ=7�2��-��{�I�Ty{:d8�g�v��U@^ʳ���2��or��{�zY
ݤP���G]�e�2BvX���!��B�*�ؤ /�j��%��r���NsO�q�,�5c�d�jaK� I���g�\��I���ެ�V��~��]-���Vì$�9�4�tN�����A�Tm�|�y��Կ��k�k����)�|}Kdܽ������ -��9Q�ܰǻv���׾V^�c������_�o}��/�Ps��"�.�}h�C�D�fȐ�������g�� �jW�3_k|�(�T�:+��m|��[@amEj�*�	�c�"��i��^{�.�d�:�U诿����Mɤ�U� �4u��B[~{ '`���ׁY攫�:08��+}۝��r,�0�9�ԩ��3��� �L����sֽ�'~�DÇ��ΙW�=��XI���ॆ���x��pPT�֮I�m{�2u�(0��`mg
�YKS����~�Ƈ�-�S�n��V�^�V���+`����XR]l�.[��VJ����^m�5��^sJa|X+g�lk
�-^ZG�6o�X3{�P "ᐶ�js���)�7�WЀ �T}���H��S=�)�֡�_Q�ӧ������	}Y􄢶d �Y7`�ؠ��6�U9vD�*'*���� �6�7�Z��i��H��S�o{n{�(�*^��1AxQfF�_��Dz�Ձ���ج�&W��Ԁ���U��Y�5#���]��<��]�ib˧�6Y������IB����vx?�4ZY�lϵ�o�v��?�x�ʑ;��=�ȅ6 �?��"&�]m��W��E�L�R�O^+$������\�Е˿)��MAU��:~����bDV�ym��*#7؃��C�y�v�G��Sme�"�o���}����f���{G}�+Y����/5]So�f��@�S������������x�;����Ŭ c =����[қ�������z�w�'��O+�\^�W!�>23�ȧ	{�{��Z��z��Q%�0�Q��ޱe��,�05�/��/��_|��K_zz����1��p��"����hƴL1�t-B2�f�0SY�)�Jʴ(�a����G�P�4�"���m�q����% �<r�[���b�D �*� PK�,Q��{��i|�c0g��ee�/[ƺ��mV�4;�W͈�AL�Ș|V���Ҡ����N]S��1�4;�eVP�!̴��ǰ6SS>�E>���� �^����{$�����mk#��ʽ,Jmk��j�5?�%�G�l�6(��K��-��73���b\u�	���'N���1+�DcV��B�Fz�.��g��낼{3�����Q����U��d�Lq2kH�@鱴��z���q��/j� ӻ�F6~c�P �?�H!ն����=��Nz��9qm<�'S�%t�hzW{	@[�˂�y�E�?�,���d|=Ϡ˾��1H�+���<��ޯ�c����e�Y +m�ߕ1Í��L)逛�K���h3�]cd�G��V�Ѧ�^�^9�<��ܑɳ����;,�^���T�K��^.l���R���ז���2)_�<���3Ea��K/�\�����~��(8�z�dB�X�v	����2p����wb��oL5�1t��{�[^�|��Yn��`7l����#�lFc��2�?�S�>\SAK�m�`������S��]:����I�� ���+aU�X��$4����2��ϧ[e?�}mT��~�׆_��_������9<���?0"ȸ���ͦ�j��a��]ÓO>9<��/��3>r�|b���wj`���6o�n>>f�/�=��y��1�n��f��=��ky�EK�I�7+�N�I�h-A����~F��;�!�a ��0M�u��U����2&�7˕�� Yؤw�|�}0�	���ݣ��ktLɊ�$�Z{�{�bss�9ҶJ���[zmµ�/:QU�`Q/����,�>0~p����"�9c�ݶ�S}U�ѻڟF�r�)'7#����f`ڌrb�;WW<RV$�M��$����W�#��\$z�I��YtBiR�ާ@�JOʀ��I�x
�R�@!�u�Ɵ�T@;�R�P^֧�Xi d����Zmr�}V.�|���T�^�k�C�S����#�K9�����Kmu�U�ncO#/��8����;��� "3�
�;�%,]���oʤ��e��];��]���X�I{�A������L��9r#){��m�s�&�m����4�uLN��o����5�oF��ɟ�+��1��J�0��j�\�^�=���?�����{�W=eʒ����_|��Z�i��6z�v` �cnۢ_�*-^����_��gG1`#��:Uh��rY`�� ���'���q�h�.�<R�O�ܢmH-��q�]���0	5k���hq]~D�%Bx3|�ݹ�,��,��N��xW� �-�ΐ�[f����m�M��T4$��'7+�V�|n�+*|�ɕ�V�Lo��k[b�@8������i%����c�l��a)�Zȑc}v���S�8�Dc��EL��&ta�������G����\h@؊ӓ�@�ϼ�)�ݬ m�Z�'7�r����.wՉ���Φ|�����xXs� tuu;�V?���GkP�ر骞���F��l��Z�.q�ڰ����M�ѯ�s�ja`O��Q���� ���^�����+��x0mq9���){m(�r������d�	&����1���WY����Ω�b� (
�e�?�$��-aP��׻�}B�)�'�z0�SMÕ�KhV&M�X�5\�5AZ�aRؚB��z����z�d9��8�uݒ���#(o��Wϒ�����椒���i"��DJ�Q�p���2�l����8�C� `���O���U��S&J�䉓u�v'��N��dK�L��,m�]FEFY��)�/ԫ|���̡�C���	�H�20�X�s�p�P�m�g�K���Ѽ�}�f��������_��_�)���<� �Fɷʕ����x��E�͂����H�}��`�e��7��@��\I�m��1�y DƊ�f�(;��ɘ����?/�G؉0I�
��7�w�xY�!�w�y�v��Ͱ�R�Mm�4�!����z���D ��}�$1�դ
��|�����OP�P&�`t! j��p޵[�����{��Z�ĸ��������oغ��rUu��X��� �-&���v�>7��\�[B�kfC�P�� �++7�SS�:ӄ�,�r)\k�
+߼yB�f���s"�f,\Jz7�{8���OO"���U��׶��?3�̌*O���H���8�z�t�V���&_y�\��)r�r����尾��}��xoo�>%���o�z>-��jشL��]V�)d��{_zgGkƒ����ѭ�S�h��
'�� ������ӮW~�z�P@w�3 Fq(gY^�]Vlh���0�U��t�C%D�z���c皉��'����C���b ���ўN�Ii띩7�ʘK�H�
��t+���a� �Ф��L����vEݼ��R�3
�����'��P�v]Z��-*'�×�q���zF�U����s���!�e�Ϸ��@�c�!�7yi���І�˅ȔM�I�ڜ>ֳ�(?}�=�ߔ?�����Ž�
F_<�2O�GB��(L��f7�9)���٬6���^��ɹr�1e+zj��_���6Y��&�����U7ȉ�z;���7J~���V�����!�+��S`c�V�R������瞯�`�f+�h�P�r��X^�������g��Y�E�D�υ��g4�)�ݏ�?,#}K��t})B��m�	�P>%y��WX]}�``V�4����׹h^V෿��ڳzf�tO�u骕+˲�Z�~�M��e���*��ʆ/�>_п{g�ylM��{i^��������Z�1���N�]c� ��	�:bH`\ܘ��R�)G1p���#  K�?N�K������/��^ǧ7o++�O�_h�mV��(LʇX��40�>7�ep�� ����v~17�T��=�XI%Z�J���X���\����/����c��3-_�6�Q��w3 X�m�� �٢Q��Q�x[kq�5��5;|q����,�+��o�oO��^Cs�]L�\[�\
�ఄ���ŏ��勗�7��< 'Kһ$@�������֬��(���X��)#�P����?��׮�v_�<S����r��Q��ܬrʿ�乒��-	y���;�@�Q���$IaTO"�PO�]ُ�)��x�"yZл�.��,�� ���v��n�G��!=�<��#e������'�iɎ6ϟC�6�D=M�`�P�mpw��	z��x��꘲�R>e�S�Z�c�V�0�S� �m���'�ӋҤ����{o�ܪC���0�s��G�g�x(�B�7����sf&ڢ3`�57k���81���X���_���Z[�l��|x��,=���������s$�\J����&�k)	�����0@��Q9�)�\�Y5������ �Bq��b�uQ�?AR�mge��t%�����G���گ����j�\�e��m�&�ja�q����"��i����#�W��O���+��J��,,N ���vzcbh�uedV��=��@tCO��qк,�0�ܹ��H,���_���0���7,`h����&V���77�n.���(�]�f�yT~�X&Z��m��%,�5������p��=�R��� �
�>�=']S3�G502��?u�LA�PhR��Z9Wn�3W��^ ^���� ��.�
yVh��XW, ?
+}��ځ��q�]�Ƨ��P{����C�Lx?�l��<W�t�X�-`���}	2�" ��S�R��b���W�?�j���/��PY��]��H��nC
���= ���EP�U�����`���ߕ�H�6_�����X�=�:�P��:�G�i
�F� �k�B:��i�s�����x@ǚ�@Ɣ/�(3:2:�:��r��2b�6�
^��)��]�~7�W>��J��7��~��Ѭ�2G����^C�ff͙Sg#'b�~Xmd]�oD�ܹ��G�Y٫�f=��C�f�YW�z�����3j��+��RX�D��~�~a�O���T��_�հ7�����W~q�������e���fU�րu�Zb#}cn�� 4N��4&³������a0Y~j@={��ܹ��|�=��%�}�[��Y�����rV�=���ʝ$?�>�h�#%ݕn���;�1|�����:3{b�V�#��Š\,��WY���4��_~�}��Z �{L`3(�g����L��Q�V�ߴ�h��~�sK���
�@]��V�Ύ��2 l^?�� ��+vo�N״F 
��G3=t��,�	��#(�T�|&�	ĕ���O.�ϼ)aL����ɔN���7�#ef�`��T��f�,>�qmX�dQ�h�2&M>~����Q\�I��6/�2�����/�Ch����G��9��)Ǵ���'O"���BOmq.����G�oݲ�zI�s�R��m覻L�k1��$0܁z�׮�1���6(.׹{�S���Ʌ��/����k&�t�J�A�
M�z ��}���W�
�U�P3cBst��5Y�禘�)y.������N�(s3B�EM� |��V�ͅ�1�]�WR��0�~�-8T�%tc�S�dQϒ�����r[�\�B&���gU)����|n?&_���aD*wߐQ)�4�#�;/E
�����q��ŗ�nL�Fs� ���8&���������c|no2�r z.�2:ڇkEdoY=�ƓV�u$�S[1,-�1�hݺ;jl�����o��/�mݹ(On�'c��R��G���ԙ��W�㙏>���[����?��?�e$�M-�Տڒ��3X��$x�1jo�����aLO(���rg����7��k��hL��<m�b�$�k�)!H�Rm��D��q��_Ma&u���������?�o�Nٗ�YR�L8�FԸ��.>�̞=o�+Zc_�u�=���T6Uη�y��������f�r�������Y����F0c]_�O�єN���\���޷j�(��˗��Fe��_�{�ۅ�L!��ի�f�^�+ٷ�էSL4cP����_�{�����/���.�q礋��77��|�{��/7�\.� �-�H0w����W,�̌���p��X�\\G?�4t�c8��P/r��Jx#�zzI��1�V�1�'�x������VM"���gЊ0Q��������i��QĬ4�&ޱ�ǒy�\��;�Wiz��kq����q�Pv�u�X���כ,�Ic��n,�4��Enl�����vl*�d+�FK�ڿh���%��YIbFIM�4E�'fN>�0Rvi Wet��e�%�ߣ� ��(P�_��� L�n*�-YȦi�v�UV~�rӥl1)����А��[Dg@�[�hi��������ơ��	�I�u%W�}�1-�t�@��`,���B��k���RH�S4��T�!����-C1�A9������_� چ�ӫ�Wz��>�n�>T��Lۤ8��='�.=�O��Sc��AY
7��չ�_��W�A8��u�th1���Mד��U̳u�~ާ��y�{���Ӱ��M�k{iԵ�5k�Ґo5T�p#�T׿��iV�������>3j3�Q�6��I: �5z��Ō�ܓ6�b[T���oma�F^T3�j'Ƽ_>��	�f�J�$���E(�EVr�UG9�?���Q|�wXfqW���q��/���HԻ�v9��s���":�5���� +�D{�J~\_�*�v�]c�5Fo=�`F�BΕC�яBÌ�D��n�1I-n�e�wM�4�(ۧ)���=0�c�T�_4��".�s=���}�����k���aL!i]o���k�i�[)���x	������K���!����j���-�\��9�	�$DW�+�f�#OZf�2�kB��(�WvY���#��*��4(+ ���+�L����Z7��n���^�}�k�k����z�+f=`Ţ&ߵ�D�ɏ�(���'�|���/�L�*VN�)���e����l�L�	5�Yp�sd��!�ϝ�^�:�?��sm��ݓg�dh;���O�Gw�?��j�zV�r.�6x��ނ�j!�:%My���fR);�ի�N^��(+��_��9��oTO&�lz�Ն����T,}�<Y$f�Q��Gʣ]Ս��ǕxA(�R����Ë������ܔ<��qm3�}�):n�����r�]�|���a�XoIz�6 gA�Hmuh'"O���]+�g��D�ͱ�b�rM��mZ�4m$F�#���n�7��ӆʁ�Kq�A-׋շ3��#�F�o�'Ë/�\@d�W�|p��l��Vҟ�Qf(��,�9��#aR��ۓC%�
ɫ��8�1tn��o^O�,3����<l޴~���]�p	X��-[^n�C��uD���@�8{����}�w�qᜋ%��	��8,�w�{���˖�Ƚ(*��B{_?�@0�sav4�r��-۶��.��K�/�������L� (J�� ,��O�H/��7sB7�^OW~�A`���q��
И��et��ٔ�'.}�B �,W���������i+�%&Ov��=|�O ?�����+D�̽ӿS��X���𤱋�kהP����GfMO��D�I�A ��	 
�A�x����|�\[��[�%�������7�'��� ��oc:�J�[���k׭-����MH[�
H��{ ~ Z.��K.�\],T�#�ĥW`�j��m�$V���K~��.M>q>E������0�6��u��s45(�l"z���<�H9R��d�iY�)��\�<�ƛ����Q�M`hV�Rh),i�� <%j��qC���3i@�E��1� _Z����w������1�*K��
Rȡ������+cx|�!�⡔��������~�_���7n!�[o�=���뛹5��Y䭐,�fѺ�e�^p��|Ǫ��|�-}�b��9���i��/�ЬG`U��u�vW%�ʞ�Ғycr�R�Ύk֬���?��?| ����c'>������Z �Z��s�ܼe�q3��Q�;���0-����&�z����Ü�ӆ�w��X�:�����lg���._�Z�d|}����a�0��X�$Q��zg��o��^�z ��������+�����/���z �G���%D��gΞ�U�lؼu�b銲���X�M�n+w�9�=2�	��/]���گ�uc���<k��Z�dv T��op��=��"Ԉ׀���Z=DE��F:� ��4:��[�1���pY%���f�0_���C=�9)�S���v���Q�Q��>.K q�s�d�mF��K%4���;@����J���m �-}���`\�PW�2^�x��R@+�7=��^&�Q9�
���]E
�r��t$��m|�M�Ipw��ԕ��R�.W+�u������b�6Ynn��~�:��<�W�<��(t���-��JʯWx1���n��1��v��zk����~�͜��z����G��ZdÆz��S5�Z����"�X圧A��l���NE��Ul^�6�:��xU1�KS!�Fl��="�`\�y;2z�L���u��[o�u��_��__����E����qt�0��A�Sce��dT�Ƃ��������x�Y�?J ���f;'8�0��T�����ã�>2<���ê���j�o|��,4����5<#L1;B3c��!�N���i��7x[��r@�P�R�D6+p�Kߤ��sf�2�?,I�7g�0+�53���X�#�עe�<p�����^��1�%������i���m�����YW�O�,kf��% �j�R�Vu9	��P������?r��YX����aK@��%�d�b����H�X��{�>>V��;�2s���<��e���)� ��ī�r�,7#�WkM��+�>?0��L8-�Ѷ7o��qc�&�=�𣥀��j!@f��a� �=� $pncBx���k�fo�ߔם1Φ,V�����	�r�W*m�����h�x:��������� ���rӔ\`J,r�}=/�R }�����[h@�C�?K��U��ʡ��r�������� b��E8�����>����o��$�d������x�*W3R��atZ���zV�F}`�25��P���l�Ƶb ����,���(��#��mՄ������S��G=�!kݏAY���XP�K�{�u�QZ �c�~>q}Tʝ.=v��{x=����:k�W�F��o���ϵJ+ϩm�y���跬l|�׆���s��j���(3�
z�5D�h|�5+Az���x8�_��s�ޓn���瘰
[�Q>�R�+c^B5�xMP>�DG$оĠ��9��?��ã�<ƷC޳�b�^8R��TJ�����r���q3̇>� ]��z�j(�
 �[�(7w���r����u�o6��O�p8w�d��F@�*�8+�|�4L�q�����7�,�v������jO���ܙRF�Yk���+��x.��/��h^+�C�z>���(�s)`�ꢕY�mÆ�5����/����P�;w�(p)�Lj��KWj&�6X�xI��w�}���gX�b��K_��p0��e�`qS��XZ�:zQ��Ol��)��&� @�j�I�ڬJ<a����Z2Ԧu��5����,��Xm4]]SO���Q��A-X��3��e�ݵm�p������4�i�,l.���o���^T����5H�x��r�$:J��c�!��00�0�
��0`���+�;%�	��y�D�p[|V=败  �a��'���@��ԏ����"�hƵ���V&����VϤY���j�t��u�ϵL-�t�W���E��n�_J](b	�C���nq�'���6_~bʐU�
����R���H�`������� ��W.��K��M�ـ��ɟB?/��#u:nt|���z;5�}sY{�_����=N�?�bD�v�gSxx���<#�+nSZQ{�V�"��%�4N��Lc�>�ѧ���Ҙi�w�n���hQ�5a��?�H[�L�1j�x�o�{��h9�k8��5�1�56�A~�'�x<���>k���Fd@�b"�5�"�\�i�)9:��){k��ҥ��]3'��=�⪹���ٙ��u1�o[��i�ˍ�T�=��1{(c���l`ڛ�J�����\@����y>
(e����@���R�yK��.S�ldWSH��}��
�S�$�^Ъ�׃��\at�M�>S�gS�O.\�zU'4Aw�J�X������4�y����7��i�In�
��p_m.�گ(�������H��I��3gڳ6��yׁ��qX�Z��vr�i�-�@��~5�5��Cxh�<��Ӕ~ 4��tc��\�뿻���X�}�f�#�-ڇn�Z֦k,Y�������\�z)�����Z�'��:�j�2�+ڸkE�I�<�3��u�on|���3�(�� Ge�0�\���{���9�[���nҤX(0�{O���ȅF�wY�z�,�R��Cz�wm���Ϯ��-:���� �A����ܰ�ڥ��%e/9W���� ����D�q�j/r��C	�+ksjh�����(on2�[�F���(C���-��\��i�@�uo��4����ڽ�͟W � ��on�T0 m*ߧ�GnB�+�)�Z\�؄^㋺K�g���A7m��d�om��ИER1Z]4@i�kϻP���H�R,���)�M)-��-��_��_-!�M]����b�0:�f:!�UWy�29/E���BJ����@P�t�<��	9�f�X�W�?Ld��F�̯W���X���+���lM���AW����哶��Ǚ3�Rv=��e�zoV��Oy�fY \��TCL_{�$г��-z�7�I(X��ŀ���S�xπ�kk֭.^XV��Nȇoٻ��|̀Š�ʔ�l	TLE��˽�vn�9
m2.Z�X[A�������k3���ޑ.K�F�A�[(N*���@�uL��Y�g�'X���U���U��v˹k��f������'O�$�~ϳ��<:3�x�&�Ú�rڒUw=�Ή�@�;���I���vmjh�� ){_�r&����
-z�xB�*���nccϽ�x��~�R��������%/i��f����)����G��T��<[���OTL�y��E�=i{)��������k׬�^u�9�)�G�6M��]�5��m���7c�2Cj^�Q1�׬��#z�>a�<��V�JL���瞥|*�*��G}�Kw�@a۾m�p�]w�0[vlC�+�}��4�_��i��b���W�����{/�'V3��鶳�6�[�ݾȩ�+�CqT ��(��gKP�I���U��Ȓ4��4:��z[=[�eƊ=y��*�|о+�YB���c:��!�bq]�|l1��u-�S~c�$R�U�Z	�t1�5h��n�U�-@ ԫR}W��X뺰wܱvؘ��7h�$nY�
�70�N���d(�uw�+����x���<O	������ j�@n�[<8�:�[��>P4w!� p��g�W�UP\��ƝDI����p@�MЮ�d۳"��r4~�0һ8�/�)�vl
?�� � *�Uv
N���4���~ J�=M�!���sQ�,��r_pOA��p�)�I�BO���pp�  E	�}(��k����V6颛{��^&��I[*�|��Y���:��ɃͿ(�>uT .xVڕ�����=�n���x�Q^J��~� *�4�n�MƔy�u�㹐d��eR�<ʫ[��0�"y�}��ڒ�Pg3�Кە��hx{�ʓz���Fp@��SGz.v�k���t��r���Vǖ�<�_�OlFp�eX�;�8�ޅ��{nkFEm}`'E4���մ��Rq�D��>h�φ~-Nz��$?�����qtwZԥ��ڱ��g�kݿ�^i�b�b�н��4bSB�|#��@��J|vl�2�x��,�g�x?QZ�Ym]�C�\����v�_�3a���?�T�-�,̫lf�, �Ƭf����+=����E��[�Xq� Ӟ����|�?�P]�w\D�E�>�EK��%�ƾVEqp�8�����}��+\�ޒ���)ĭ���c��;��W��\�����O�B��Y�и|���Eii�G�o�o�����
 �,7��W�6��g�[\ׄ��(�v=��������5@�f�ʻ���6���T_6E\����(������?B���X�����;��ƴ�[�7<ju��P�$��L��m����;H[˷�'O�)��6`���ݥ]����f)�Km��2�R/���E|�
��9�-�zUF���u�i�SoG���ձ'�����я|���=���}�W�h7��~�Y`��Ҧ|?���]����1�ZC ���D����p����]��$Xw�N�UΦ�[[�6�m=��2��YǦ@z�{l�Ԣ4D�$��{���
��l-
h7���������ތ����@j��㟄%$x5jU.��E��J���f�gD�;
�`=z��Wމ��*�2T������
c����,e�<��Iˡ}��`ͷ������[��e��v�w�/�41eԊ�X¢�����^�����-S���}�VI������'â��ƍ�zk"TG��z�� ���f���8:Q���}���r ���'�>�hgO�x��ju��i��w�adf�ݦ����Y�m�Ϝ���&�a ?����{���WU
ٖMa�&�B�3��.����p#���-���^G��0%�'���\��m;g� �{�<>%㛬���Q�|�Q�D�m���ђ!YG�D5|�Z@�rhx�f]�[��,i��D��n�G���ʅ������fVy�- g��A����&4֡���[o�>��w���rM/Wv��Z��N@���\���Qs�m:�Y���kNV���(u����=JOM�T�s]9(y>e��2�x�"f<���f�{W�{�a�K1�Vr�z�zJ��Ak�V�\V�ӳ���悢g��6U�.t��iI_o��d蕬Yn�Դg�C����|)��)ߦ \g�������}��u�7�Z���[;��X���ڞ7���z��E���QpM(z����.��ix��ӯyGpM�t��-�S�%*�:	�?|!���槟�����S�h���ʻ*%� ��K&T���g��XHzE���D\�>z���wˢ�ؔ�����7�{f����w�}�<XS�̏�r��vI�� ܴu+S�B+�hiȳ�7%�X]F��Duu�B5��@+����t�őˁ?���˦��Q��.�(eSwit��ӵM�1`�۲��ʺ	����m^��p/��_>�ܱ޾KK�2W.����Z���$,�p�*�׋08ج}�6h�>Y�Mx����vTv����h��@�:hB�nqΥ�W)Zuc�k�Χ<3��9umL���-]�E0� 𬞜�"�׾G�B{+��K���)m]\[�Mb�D�g�V���hJ��Bs�:񷲐%J�v*[�n-E�'o,~���'���d�<�@~��ؿ�x`��ڶ�w���|���� l<�V�Rƹ�[�p� �ܮJ��[�%�[5�y�%
��'e_��<+}�V�&}��@�Oʹ^<��Lү��sڅE/��U��n�:60>�kxBZM�FwL��zHc�J;1$��aeWh�J1Q��O+��z"��R8�W#Џ��94�u��&/��םw�	��9q|���=�_�*W���d��(/��Rv����O��i2X�e:^mp�`�-h�t�F1{�+�a���U�4\�ѳ%8U�	�d�Z�˿���*�0be��*W�0�2J���ʹ�c�p���(��k�o���3��0Ȼ��ӱ�����ny�1��{ʠqz��l� mh�O�]cU�X�v�40˪`5��6I��
�@=G3I�ϧ�_nV7���ô]h奀�W�>�X�w��i���X���e��#k5
#'暑�Ј� @=�6_3:6�� ���L=*�}}jQQ�@xc�}�U�ĢsNK�C����x��v(���K����\�G]�Ƃv򻗷�3el��Z�fehQ]�~�7r:�W2i��\����'���ُ�Ն6	3;i��58��z��}�d�;7o���e1�� �>a���2����}���'M=����]D���K�z��&�c����}���M�?��E��3�8�GG��G��g��������#>�����S��=�lp�᧎n);^�%cn�ڲ<
So�q�-������B�VFh0��d�4�����8�-��=�n3<�����娇�ԥhExot�LҮY=����6Mz����Svv�{�;]�(K�X�p]�%0c� ��:�������r�-&����Z��s)A��O�Mw��J
P��T�">��:�+egASd�ֳ�o��#�4�^�#G��as�(W�k���y+#M=i���i���$|�+m����(�kW[=���@��{K��6� �{@�r�Jɫ����Z��M̮T׷Y섢Տp��众Ӕ1Gϩ�|���ѭ��F�S�j�7	ڂc���g�I	yh��ҙ�)�X/%�#@Կ��}�x�ȝ��FA;v�O�I���g��;����{,c�מ/�J}�Aw����W���M;���D���V�!a2Ӊ��S'��@v�H��*c�e+h���k
�����a�:�[o���R�[�M�7ծ����a�(��,w���%���|�$Aݫ=���~����S-���V]\�u�]��и?�бG��������
ޕ����zϻx��6c+ g���u���U��rDF����!U����T��t�To�,��k���y�)=�Z��.����h״o/��5Ɠr�VY���A�/��������#�t�����:-�"6��x�#>*<�{�i �î(0f�5߷�0��B��{��rh�j�"��k N׽�rZ�eT���s�y���y1�J�qJd��{T��Ⱥ���Dҵ�L��vfubv����l_�W^y�����k������e�,K*B7b+O�sZ��/&I��-�4JH�F�w��~���?4K���$і�f�I1:��@BDk�n�@0Z4����XT�s�z)��V�ǿ����_z��S��uL,�/y�&�n��VP����W{�Yw�R��-�ZFO �NS��|���Ε7�߱��@U�<7Am%�|�
P��M	�&]�%�KM���)�
�6[	�ֽ�F>��N�òf�M{�Ѫ�gs��PE�G� ���둀~o�B�	9�	>e�v���fh���5�a���1��[R>=
�b;�r�b�}{kl�,"./���ET�2>B��Ե���X7�r�M`@�rwzjea�xǽ��g�R���#]�u/�;�� �[~�o�)|.���*hk��"���X��ԃ�`>rd��`y���l����ƪ�DA�G�7�H�E�'�mM6��s�ֳ�U�Z{N��v����Nu��M������W#Mm�h:w�Q�{����y��&���q1��}a�g��n�f��m�|�ӽ���j�����1(cp�, d*���\�e1��q�۽b�~�����	�jUx�s�[q���,L���裏_z�K�C=\�X|v���}�6���C��̮iZ��ixej	�V!vc�iS7&l`\��`b�q���`�7��x��m�����͢f�����kK�"6�Ʌb `�f#4&��E��WY�uӄ�1{zN��� fk�ol���LM�]/��3��&�1�v��r��}�] %y�0m�$'�\��ȷ]k�W+6P�<��ޯ�*����U�I�+�&,�ꮗ՘��W*�1����x�<�6����h0�wշ�O(�j��a�{s�t-P�9����W�p S�r����yт�z�z
�U��Z���2���"L{Ԗ�Q4)EM��4B�~��qA��_�R�j7�y�����g�U��.=�W��$OK��(t���G�����	]\S�j�j����(����J'�[y��>c�tt���x����������;������f_��\m��J����d��ig��p�f�^r�m����M�7��+\�f�->�d�gam���`��O�i��׿^iX�!��_m��-ħ��^�����o��f�tC��駿8<�����1�j��ɕ�0G��\��������g��k�R���y��� ��Y�%��_�-o���ͳ�O�<U\���kfF��5����5�|s4�� �+��i]�O�(�WV_�#wK���3�Ϋ��^"�g�E�R�U�����������BI- {k/= �{�����.e!���{/mf�h�'=���K �R�!1L�4�05A-�*��PB�g�m�wկ�i�T��>%1�ޘ6+�ʿ�!gEO�O�G�\�����z�?Uq上-5��1��;\�o�a=���ׅ�c��AR���R�	��u��Ғ�X>�B��3~.(Z�o|NɛQ z�Q�I��c	st�'�}�b�ɛy���qa"c΀d}$FQ�[���H�� ~�6l,W��>)c
�I6Q�{���B3*�_��(���k�h�	tl2֬�R,��vo|�4�rV�W�G�Ƨxy��%��]��~-^
����깑w=��.���r���?�_R�{Mfz~�̣�vz����o�3@MM޽kw}�fs�l&0�k��]G~yԷ,�Т���-Y7��P��*�RGu��<%k�?:��������k�S_|2m���?����V�T�0��h,��|f��Y{���U����>fɰ�3�Ra��(��#0H��b
=۵0�v�)�iﴆH�u7Ybxو~���v~����G��|�s۶T��^�Y��/�N��S[:L� �X�P����{�;���1�����D:����.�ť������|����{]�d)�ͳ
��|��t�9b�A)��JQ~B@�X�B��őY��h-u��(����]Ϥ�uT��K���Ő@���]�r��<��K�fS�ؒw�/i�v�Z^���ϟПq���8���:s��=�*s{t�|��c�z�S_�Ԭb@�I<fV��c!ϴ�Ǟa�֍&�Dq"TF�� �v�=���da�7������z4.�-c���95k�k�%�z�s����}�E����k[X�����uZ56����\Ax�20^���=F�g� ��6K��F/w�{#_y��g��F�v���P�QDi�T�G����'��q�=�n�o�_�q� h����x�+��L�e��J;��Js,�����.�;�[{{�`5���]bMS./J^jn��~�5�L^C���-}�M��b_0A��D�(�|������|O��/��W�/~�r��ڃ! ��eǎ��4�= �Ȧ�$둕j����
��o������(p�%�kǎڶԱ���t5BQ%{�;�UT%R;��X�#GLV
�����mٴ��c=�����ݻkP��8p���Z�4>.lN8F,�i~[�)��'�)��x�� 7�Ntmd��D��t�6��$j 
P�͖���×���4�/_x�a۝[��f�؊��y1<�<([�UV2c^��5�V	V�=��-F�Kq��e����^�ƈI7��ݬ�&�_EiGx�m�iB�����F�Mq������-_N�tk 8�B��[A+�z&�$�c@�2��3��8�U�F0��膮��z5�F,��h�6�=�ËT��5>�A�Z�ƠX��s��zT==�Z �̱&���W6ͳ��L�ֻ��ɦ�
�@+=\.���mz-�r�1J�b�#G��:�I�sm
�z�
aejFa[��L�E/�W��(�j���|W�4����w�yVP�)Ѻ�^�g��u�P����_�D)W�~�ѵyn_y{Ԋ����[ٚRj�n���	K�s)sz��Cl�'q��.V9}����^y��2�)QrͥFqnH4�YOD(����)�ŀ���)1��?����RJ��<0�nc���Ka�L�hi���|޶-�ܜf���K�k�o6�[���P�92&7� {�����g�o�r8?,Yܾ�˽b�<�h�J[#!ZsgX�t��N�� �oB��%@� +q�5�y˖�R����j��U���?�{��~���|���lbQںtiF�!Z���+��1�ܒ�`o��l���%�j�@�iY�	:��v����>�h'Nۿ�5,�����g˰���[���W�Q��㷝�C\K�����ӦC��hC�����V��й\:y��?�yu�S&4�˧�iK���y������gz�ԟ:Q�JE4k�+y��P�-��� 4[#��E�ϔ_�@��+y���C��W�1��t+�\�c��1�JYk!��?i�Y�۩��z���[�F;��U:w>�v Xʍ6����DWS~*�����g&�������q�9�Q�*}~��_ƒ�����z��4�o�]TӃ��V���ȍsys�}S�D	Ɨr�.m=�RQ*��k��g��P=��e�m�Ԣ0��2+e/pM, �5y����b�����~ZC�Ƈ#�d~�m�t]�������׵%ʭ�yN�㕫����5V��� C��f��������H�m$��s�fSI��x�l�xs��f�n��.W��)���\�������/�<����W^zq�p��p��e����1lڰnX����+�/�8
z�����	mP8}���-�q���ɒ�1�N�KV��k~�p��u���Ǜ�?|���=|��/g.^v���p0zպ��;1���?�?>�Xk�9s����A˿��4Dx���8^�p�����'ca  �Y���.��Jf�FK�E��7��TT#��V��I��F���"7�Ծ��v����{wGkm�Q�-[�,�$ z!����������_�s�ͦ/�~���N��~1>]hWI�
��3@�>ט�)D1�D?r[�ee�6M�[�`�7��.(�N:��#F�)�5kקW4+�;S���{Ӓ�ǡ��+Vkô��.�1mS<;����ҵ?q�x�r�|vv$:a5�s�Rڕ��y�>Xn�����z՚�{Bĸ��e]Pm�������u�e�\6%����b]ִ��m�YmM��C�8|ٟ�۞6[�2Z��C,mm��P{������I�jҙ[;�~p�{��aF~O� \����6�n�hZ��S���'O�5{��h�b	'���������k''@�~�r94������G ?"�F�.=HJ M�~W �L��bBｊ��r��1���j�"c��o�Ў�>�h�hIڎ��1�a�/��,�Tm���D�5�c�JsYޗ�<�⻡z�����}� q�k��F���cJ��sMɅFN�)��5�m������j�06 �6!�G��w��ޱ-�'W�Ӂp�m^�Gw��6/�4�sgDF�1n�ޱ>2�n�Yݚuw��]_Y1��b��-��8W�YWJdy4qY�-Y�"���;�X������qU,�;V��G���}8�͙=3����[M�&yq����Y�L[_i�~� <�J�fT\Ϲugk[۝�m8Iv�G	ز�G�x��85������»7��V����t�����px�W����g�̞� L���jՕ���ـΦ ���Uِ�~S��H�\�׀��	Cj`g?��T�UaH�
0̶�b�z��3~Di�o컩�פĤ�u���ٳ!ԙ�g˗y�̹��Z]��b�11��BuQs��e��oV�D�Ƶ�]+��'+��@
�K�X�$���c�t�w���N*E�X1��?�A�7��>^
bQ�qg�V.K�+=�Ea(z%��[ ��ُ���Q�Z�/
H t2V�"�i@[= H5�ĸ
�����.V0�;��Ȅ�	��`�_����D�AE�S{k%/^2ACt� �����׳�7m����u?}���s�&�x����w�����C}j2m{M�'�I���-~�	�c!�\�[;A��á(/n-��=W��ԅ2 $���v4��8�x�Eg�C���ň(C��$�v�/�5��A;�O���(�ozN�/�H���r��.�����( ������~a��e�C�{����932��Ѝ6
@]D 4a��=�;w����gE<��T9E_φ��}�L�Q�v��K�\J�{�kE�Фʝw��E��[�s���&ހ=k����	�G�zq�'.�;���0ch���e���ĕ�+V����R{���r�&-��a��������;�6�G�.�7G�R�'�|���vl�6�]wy0i�V�oV{�k��U&�YF�D��f̙�b�o�hl\R���|���W�\���������s��Μ�0��s>��I�9�k������B5;���SX^>)�2	mٺ}�v��a�Rٵ!HӒ���_8�	�!0ȪX�x�0/�][kpI
V�����b^�۱R̓$���Y� ߪD o��s{�o��ٺeK��;�YX@��]`̥��]�~ݰk���Y��KcZ�j�cY�`,ce��4�/��S�,�s�2�d�Fj�}bF�g=t��w]������S�<
�1B��u�}�eo�Z>B�iae4��U+�����.^���H���\'�??�
�ة��[��i��PZ��x�z�Y�7�gz�j?K�1��9�
�.b���Nm�@p�@"ĺ�/��b�R���#0,�U�)����EbL�����a���_=@J�L{i�)���i�-�=y�t}m_z���\/�-R���p�Q���2(# ch��Y�N��.��m��`M�  �^��!�l(�/WGz�H��h%����&���i���R�+#��1���i�����>�6�D�����\zz���z�U��*�ۘ�:�ؕQ�w3/u����s���_^�N�IsWi�^#�&���	+����
F�|�>cD9JaM���1���O.������1�����T�|��(�6Zєyw����8}7u�U�]M/S�b�	�f�vze����;�n	�5〡f��W~��z��Ў��s�:�s�C�����yO�y4|~-4�O�������`��+KY|=�K�,��,�o��(غ0�D!̋��OSN���l��x����Ji���O������y���Rpa|�ɕ!"9���/K=m8���|zp����/X\+b	�n����+�0��o�����G聺��z@�����Ji�H�®��]=��}��W�iU����5��0@�,2�+eYG��P�@{@��z���muy˚Z3ܹm{�xkR�[�۽�.�a�>���?"�L��硲�3�*а����,�?/Vºa��5�����9%�A��Y��_>�8�pA�	�������(]������C��;�)��!�x�Y�/z{�Ґ�`����E�.�4ۀ���Q<��� 8|[� ��@�'��՜�k*'w���1v`�@t=����H�Mڮ߸�>y��>���tZ��U�e�k�C�
ȡ[ە2���r�����V)Q~� #��7!/e sʞR��{�q����,�(e�'�w�@:�*@�IK^��}�3�)��U�wɘ���`Vf=[�Vb��|��|�Z�;1�C@杖Cd�!S�5yϼS��Hi"��iϠm_�(���=���6Bz�(��i�|�Q7(1�����i�d�м�����_�3��ĉS��:�O��o�~�{�P��(�I��58=�<��6�˹gN�>[V�(��������Ir�m��<���|X[�0�W����f{��A�Qxj�p���}x�����?>�v�9�>/��y\s�
�1Rӛgls	U�7uNSV4��ˀWR��)g�(���Uc1��|#5�9�o���<��"���������ǣ�ϜO��>:��wp8���p�y,���Бh�S!�'���\�Gk� �Z�.�GG,?:�y_ �üs�f�[����gS���>�O�,baj��.Y��1C�/֥����[�m��C@S��q�IT�_��sil�dn�@�(	���=?o�O*�aҽ�=���6��~t�@/f0�S ?�{K�;{Z6?�кg���הD�#c&'�+bl�NO�̩a�X<�~n@WY���`, *4J��3c�j>��|M��+0L$@@��9?��HO�ja~w�%R�'Q>zE��'� ��镗_.@ؽkW���/Y���+�	����(���z�W>��|���o�>>UJ`��5Q�_�H��Pz7�Ξ",�[uy��m�.WOD=�C;.���Φe棣�7s%����ϳ~K�8u���պ����|j] u=�"�"�*�n	&���� ����Ll`�L^5��X��D �@�߽f�]i����LѬ���W�h�9�b�yq�cS�m0��9<%=~|� M�G��צ����Ne�'*s��)��0���\��{A���/y��}�,����Z�ըT��~hw5���Q�!YO���2�B���|���.+�x��\C�S���c�M���f5��	,g
0�A}��I���!�������+z�N���M}������8|T��T)9����ڸi�p���rk��׿1�����)sz�.^����_Jo����9?���>{�)��g�^��L�z�>���RV������x�E�Z��v��k��{���w`x��{{�p�w�����w������X_��%
�?�J7�Hw4��H!��F=�°��;�s�퓎4�=۷o��Ԇ��ڲ�ر#!؞ Tۂֶ���/�8͊ж%��|���R�E��_���A������1���륝1�F�gC��)�ư��'�>�����o��^���΢-);D���W=�'y���#n&�E�f�Y#�������>9�(�l�1���.��o���W;3J�l�O뻢��`*��;�s1U���,�!4�8ڌ� ������VV��@B1�ӿbŲ�H !�M:�=@�꿏B��(�)�m]|֍���9D�Ǫ!tz'\S쎆�G��Le#����Z�b������c5#�r8�(=ˢaY3�JFw}�;��s�����Y;��N�v�z(����G��js�8i����w $�=�'_J�Y����&"`d+��C��*�)�U 1�&ֹ��5��r�͖�#�^h��3�.�������k@�oSEPJ#��"����YÑ�(FG� �:�u�<�>�¬!u/7��*l���U��:&����fx���]3�(!m������zk���M*����k���(���KYW�5.����a)3�x*��7k��dU���sa�if�9�����1cf��=��q#�y���[r����p>vA}��j��W_}ex-x�ʫ��S�M�����_���`�᯿���.�B�[ӆs�� <���SQRz�?�1Dq��/����E�T3���$�c83������ZO���"�~��0�w����G��O�:�v�p�V�`3B�X`�C8~��*b�^t#DFG.4�B���ۦp2 ���?�>�a�~�f����$`܋e���,!}��w�}њ���X~�[d?������w�q��tE/���"Ȭ,��Y5�|�=�K�^x�0��a�λ�G~��d��Wo�@���]��a�cQ\��y�cæ~��ko�5KOfђe��Z1��m�Wl$�\�Q���L�͢r� sɤ��+��X�ӻٺe�0+��Ʌh�D��p��5R>��Ǻ�m�(�Xc���Oo�+�x��>�6�f�{�0��H�����V�},�$7��;�[�4^sڲڻ���bFC`ǲ�k^�᎜_J�1�~��{�[J�p C�����}��K�⣷��[o�=�I}����\fƈ��_P%|%��n��!�MY�|��m�)�\1o�IO���c"�\�>%@V��,jn�RI�����Џ��00Cw.�Enu�L����Vȉ�j�w:xJ��i7�Y��/�Q ٔN��M��g�=����+��2)�N���U/#��6p�����Z��ª���)���'��i��7����z�K[���.hĸ�p���oƑ�]u��t��^�GI��� Е���ـ�zLyN�:��@]��'�VS��"*N�m�W�(�h���5~��hג�E.��ۚ��ۚ��$�^+��g)����⮝���}|�z����<<��K��~:�[�$��0D��1oAS<�R��ySY�N�cSx��g6�Ϝy��^"[��	�
4�
M�ෞ|x{H�����<\Μ����$��Dd�b5��4����-��uh�W�*����O�hIߜ�i�io���pÆ�ђ��bdu���,�a�r�JD�X��E��1��b���C���G�q<��p�)��ƶ�� � �zx8��;Ș������W���4b�����~W��X�o���d E�O�|H�s���2��
XM�ʭ�(��,�6>�I���c�o�xǰ}ۖa��Y�c)��x"Et8@n�D�%OX�4M���'O=�T�k�P���t)]#�+����k{�cZ&5[ �at�M��|���,D�d����˪R�|��1�
L|��٬3�.����7����ۓ��h 
0�2F��gD���d��X?�M��>�L��S3�B�`@�~��cP ~�"|f����ޒ��X�zƒ�#��S�1I�@ ��j �Ք�(�d�Y��^�j"e(L�p>XL.�aV�ԣ�����<䫽(��y�]K/���g�9���_:&4 ��t�Gcs�Ɋ�n�:�=nӲ�W�20�Ke�up��W�����zi4U�R���������k���9[ǖfʐ�( ��{5����Wh�ES��Z��
�+��2�W�U=d�k�ر��klk! +C��n��	��g��X2��%���^��Y\�(�[���5v�J�9����G��f�����O�{��_	&�(�� �0#=��
o(��Xɷ�4�^>���z�����ax��#s�$n�y���?.�?{!V���Õ��@A}$<��J�L�2r.�$5����|�!�QS+�����;��ݴiC���aŊ���O������%Q~ؤi�-i͋ ��v��;r����b%���|ه%7���'u��~������i����A�8�#,V/�4�ݻvD�|xhx�ͷ�]����Qn�={�pr��Z�����:���߄�1!Z4�M)S&u�`i�(�+���%��;kF����\�����(��|��oG9�̇Љ��`ߗ��e<��aZV�g�y��@���˱�W@�$�¬�3M� 9w��9�f�H����V,3��@��\���5m�l_겝��[��>[3�����?��5+�2%Ͷ�ؙ.�i��R2���{{����VϑPS.*h	PB���S�r��DL!���R�;Z���f�	ڮ�C8��4�6�c��_^� 2EJ���9+�*K�kJ��S|������g"Q ��=F���Ip����OS���)�~3
(ci�M�r��:�=����=�����|�Wn�q\��Zj���oc @�y��"h��G���竧�zv�_JED=8��(	�(c#ϴ�
��)w�f�P,K>�â⇼�O.��N9^uڒB
��Q�6��߰�|��f��R鴁����bF����-��e��5�i��Vo-���q��ᮻ-pM�w^�*�\�1m����Ë/�V�� @�g��M�^kVn��'�����H�p7��(�V�piZ�z.e�Dԕ�����q��a�o��?z�ȑ�Ù��Y��X噆NMh�TA4tM�J�ٸ���kZ��N�^M�ֹ^�nw�|�-޽{g �?~h�I��u�z��_0YJaǎ��X�+W�	��4���0���eZ_`�iB��o�ά!V�s���{��`�����V����o���p������o��1�5oz���~R�49�b6P�]P]NK����n*��h�A6m\��ߎaݚ��� �:<��c��|:Lb��;c,) |> ���O�R�p�����Pk��9V�����N�۶�U;/R"z���w�[X�6�Y=	���#�� �����I)
6�S�#G����x�*+�Zx�����nKy�{^3N�5�v�.K����o��ߌe����ʕ"�=�x�żd�-�ᆢ<�b����&�����Bo�4�Q��3�ڧu.Z�(u�4����P�Y��$�Y�G� � Pm�~(QJ��r�$O��6��  ����(�J
Q���4�\�Gyx�%
�z���X���4��fc���)�@Y�i�=(U̹�X5�7�p���mF��՞r�ǳ���IW�[��^�ܫ�y���&-���)L��#"&	ȷ\3���F �����FQ��+c�6�XM7)#�:I�3zj���)m�2;e����PB�a�Q;H/%�g��}�!-�z<U���T���Y��M_�.�P 8|��H���[���5�o�l��o��x(�ۆ'����Nz11,��V�*�����䭼��Vȃ?�W�Ƙ 0�p�q�0�c!os�j�W�R�������3ǎ�.^�8w�p�ҵbD]/����X��,��g9�E%#~$�}�}L-Ә^f�86��T;}g��BUP@�b�U�w�b�4l��\+p����W�an￿x�Wђь���k��7c�����+��f�?�n��W_lJ�WυO.�E{�K���o�;<�����5����>�5��,�hT��V)�W#�����D�-F�f�aN�h��Z��EM��E��\��s��� �Q:�f�ƴ��`z9���-��P�����E��-�V��O���t�Ϟ�z������m�
pÿ�<(��6�'��/�Y�&n�����1.�w1��|���f<�@5A��ݴ7��49=3�n@�,]�|��_��5�rs�P=G��Djz�2��D��|+˳�
h���@?qwlۺ��m�c�X������ܬ������V`�
d��K���<���ͩ�������,<�5�a@�iw�e,�XjbOW@�@5�U�����Mz��QN ����(��z���u�Zy�|�kE���+G`���J ��%�g��ґb��.z��{GO �^�8�'ϣ-�kږMIo�1$�2��X���@�
��ɬ��\�ŀQVS���L����L�g�H}R2�Z�4eV`^m<�Oʊ�����!C�@����n�,y~�0@~�\ۖ��-f��=9���p������%��O�>����3g��~Z���oB�5+ ��g2��)���'��6MDk��y -�G�V�7N�7�����m������/�?�I�z�ܚJԘ�5� ���!�g�K����a� 9�k�tQGHs��Z��	��@��mٲ9�i|fP�Y�s]U�T�W�˖�c.�qN�)�:�J����u�/`��z1�\sY����jᓔ��r��ҋå����*�����戛Jv��њ��Ï���Y�����D�����}kS_�T��R��&���YY�)v����TC/�j�MQf��XWBhJ(� ��ɂ�w�{��M�eQ+��%�wO��/	t�g����a��_|qX�qc���3	�>t����;{���yoxo��(�w�������'�Sr}tb���7����#�v%�����W^�|��᭷߉��V�ݻx?Q�W��j�k������\�N�ޱ��� �0�b��2��c�[1� ��՜��63�Yl�vI�E�ࡿ�h�,r�o����$�t�G��mhT���:��@#V`�'/��&a�r�iGIn
���\�%�{s�-�c�z��ZU��B�W�.�{]�|>N�l=�ܓ_�k���0���8�I� �%��]eO��k����f�O]�z�l��T��j��V4n��&/�% �Ѹ�#�jKt�ޭ �)��r����Cl� q��m�~��V3����Ֆ�����w�L�Vmg��q6?ﺯ�8#i_�v�&>Xc���g^�����~�|0��2&_y������˯�:���k��{n��/E��,y��G������"�!-�7�!2���m-�ڵ�1�ԥ�@�L�~� F��Z��`)�k��u��U�I�=`c��� ���g�h/M�Fe��i�d�Bi	.��4&�1}�:k�u�z�Ϙ1'�tu8��O֢��5U�ԙ��V����s��t��Ă<y��p$D:��J����z��O|�=����4���gN%O��k��u�mذnX�ڢ��ba%��ٽ��?lشe8K���R�K��Ƶ�Z�(?l�ԑ0�^�@c�� �2p����11����ϳ�tݯ��NO�XM�=n-Eh���z ��b��j~�w�=,���g�|��2��Q����&L��h�2���/��n/Y:�=�I��ZJtOzP~8x(�=<�07���Й�m~���}x�?XS|���kŻ������u��>c/��e�s���
s����Jc߁�Ͷ��՛1�,-�:?:r��g*g�����؄2��6н5�׀�Y�۷m�s3�����f� �����o��~�(k!(eƄI��,�����m$)�� l�/0�\(@�^������h��d�Ǔ�kν_5�|�������g���*�<��ɱZ P�P~�p�ʛ��Y�%�<S
")��>�9���h�c�&m4(�<�ȝbA�_���S��'"M��֬sQ��+�ҩ�����K;:�"ny���u�ܙE��|%x`|�>�p[���-D�r,e��p�4��i�k|����D����?>7�Ğ:��Y'>>]�r���dp��3��xz#F�ȇE������u�1��73�j걉j~[ʩ��k����myHV�ت�ì�����Fw�B�܈	�U����\�'cJ�6TIi1�1
�y�)5V���O,cV�y� 𙃜R�hn}@'���cU������r����s�'�� ������Xn>P0��T�5��&}t�}�V���2�?��ۿrX�v�����F1��m�R���d34;T˳w�>�L�+�t�8��{Ӧe�h��b���ӽ�Fn�5�#�Fj�X��o����-�)��ؚ�u���j��\�҇��}��Zo �Mo�rН,�K��<g�ݫ�0�f-^V��� ��)s�/�B�X�T��i����r�Z�掴ݧ��I~碠=ǥ�7�hj&����e���]~��g��\M�յU�Zt 0�H�kH�շϟ�O��[Q���s�%�}+�'-��,~�o�4�W��I���/۶0˳}�!+� =�����D 	����Hv��H�<��w;��5�֛���ԓa��"J��ピ�t�#�k�o�;@L���b�ɳ�P�N 7�d��H�=�(J8Pc#�[�c�����-ЉUo*'��\`�U�����u)��C��0/e���<u3_��-�����ݦ.�`�M"��M��W/��q�Rznygά���.��ݢa��c\6,_���N��K_PWJ��ԔJ�6C���"�[���Ü���jJgh��݊��dF4�jP�ծ�1&f�|��݂��N��SeG��߭[�߫�I��f�`�[�6�.<��6߼z���gl�j�k��>,��E�8U�A��*1��j ڤ^cZ��u�)	���u��D�B���������Y�,��	��?�Ѱ?�����Gc}����.ƚ4���o:ݦ��kИ�z����sgO��=wغyc@��a�λj�ؚ�+k��|��;�c�����a���k@���ިA^c��kJ04�.+�O�C@=N�%(�5-M��D���#��`,^���b�5�?x�:���ao#E	����-���{�8�%e}#
�K��={�]b�5ߡg�X��,����Y�qz�j��"!��H�Y�$����p�jK�/�����lz��(�vD"m�on�άRHk֬��\@�4���[����1U��{�2�Y���ފ*�ϕ��U�ӕ�9B�]0�)�>>�?mۀ�rs�v~}
H�l���,�f��e�����lĉ��
Kl��H�JÀ��n�z�uǛ��ϕBp>�L^���_�����GB<��5��X�Y�!�	P�_�E�)���>J��3�N6�K6 ~�]
2���:��Ƣ?v�X-�4l���%m��35����)�%Q���K9qs2:.{��v�5`�6eћ�k�2��ׂS��@�"�;֭�k[M��u�]�λ�?x�p߽����=����]w7��XS[+/[�pX�w�\6^�VD<Wo^�f�Dn�e�]�2'�aP�	P�f[�+���=���oK��N�)��opsE��p��0+�`���i�q�b㾲ˁ�D?t���m�F)��|z��0�7~�<�b ��b �6)�c}�;�"�y��''-3¦Ud��w�$3�}z���4�������"�����J�8x�t㒲H��t=b�T�z�L5������<U��z=ݮ#��Z�֜�Q��N~<�8~4Lâ�Q �kv&V��X�V��dq����e� ���)�>�Np&c�Z-�i~�r3�W�O缽c����.j��P���(��47�Yu+�}��LO��H�\hw<�>��	��^z	�,�?:Z燢DLKm��X��üU��#�˷h!L͐=�^[XH9 s-��X�d��Rr�����(�iy��ޡA��γ��W�y{���Q譙y`?�~�6���ӳ��� �p$ޫ�@��I�	5��{��,�[�n-��5�.���ږ��~w]J�Pjc�X7��,�>d�V�_�4�m�+- �H9�;�*7��]��UD��L���Ώ	u���?=�͔S/�r�'�^~�i���"���~�C���5Gה� 9�Fj�\S+}�V�f�ХL}�ݶ@�.�˗-�uv�DWm%�R���fƜJ/�TF�ȲG
J�����'�E���Z�,����}������O}ax,��߷{صc��m��27o\�xǰ%��wn.�#
`G��m�}���e��o���h�#�ǳ7�!g�RPfB��׳A������w�uW��Bz#p��Ǯ(��|r�BҺ6gX����bXs��a}�Vac�l�Y@f�b�`����6��?�௱���7���1���wn�4�B�b�%u���Z��+��L��A�`�¬Xr]�H<\QV�������n#�(�)k/V؜h��i� ]n -�o�xݡ�g�Y�l񏏸$���ʗw���� ��Gs�ư(V��y�jp�ԩ�ù3���p*�>��ӱ,N��,�K��7�.4@��4���A��KH��U��HX�yIL���\��S^��� �.��X݁�zUM2��Ĩ�<{-y؛�P �^6���� ��=��}!7���2�O�>ç�|t$��6�+S�N��I/'yR>�`?.����Ms��Ah>J�>2�������������t�2��Q�)�@�����	Y�Q+3��)�W��3?�R�u� �f=���St��]\o����0Ty���1P#ȦGʀ��Z50HI��W�<����]���W�Ɗ��1r�z��^K��f�W'���*#e>&���S��i�+6�2�(��ڧ�B�K�C�F����`v�~,l�n�FKrݢ��}����}�0	���m����t�5�M7U��
ȤZI���fU��9�7��[�Ѫ]b(�7���=kzM�~����������vﺫ���-Y4,Z0;�r�!J⶛z�Q1�X�3�֜�Ӄ��ͯ��@��<��ZS�N҃-�g�1������HQ	�>3�}���λ�js�D���_�/���䩏�o�TV�\%��p�����U+��)�^Ȏ(#��f���S��l��P���A��V)��럜3��}����<�<�`���g�����k��;�,WS�XU;�o|��B#b�%�$���~(����յ/K��G)�r4r�����t,n������9"ɪ�|��p������R�Oҥ����nY$ϰr��Θ2x�@��O� �F������>�5�&�n���S���J��c#t���=G���P�Z�6g���&k�� ��� Kb�0#BdP���j�f���1LW�� �؄$��X$�2|D��q��˲�?E��)��ź���n����;�݀sf�X����m/����BP���y5��B���T�~ &�\HZ��<��,RXy���3�k�!����uߌ��-�t��*Jm���tr�����5�1B�zU�(��?ק2��7���>UޤYe��g�s�X�!7��s=��M}�����_^ ZuN�!&@>u����0�F��|Ki�;ߎm��0�]ʁnc��f��S1.�4j3�><t��~�n2�
V��V�~)�4�WO*<�ix�����Q��V0��. �x��� =L{�ᇆ{v�*y���`��p!H�MR�I_~Е��Lri�}̭��j��ۣ8��(~�f�������bD�O.$�7\��w����8�Y�*�a��}UO��+��a>��õ�mk.� �mNV�ȾC�ԉ���s�k[w����m��6�;;'�j��5V��s�����a��OO#��{�]w���\8���;Ét�V�.��C��I���q4�����]۶Ǻ>�BjL��g��p�`�bp�F�&7 ���Ej8�(�gs��ڼ�<iM��Y���S��r72Zo�-V����Hq�4�ҥk���kVs��������g�_N��-�&�Q��e��?#��M�rꄱŚ������������$ i��Q�:��V0 �ʷ�@Q
y�#;V����Y�ea���U�9)�����)a {]����V��6��Ooq�@)j>��ad=��Y�翴 P�Q���vc�oGm�(�h&]k3�)Py��C��y����:6Z��8�=��V]Lr�����!4+Ǉ*�ݵ=�O�������}[[��(x�KFݲ- d�Ko�9p�� V�mt�*�$���H�Ś�w�d�x �&�w�t<�r�I�1�w�W�NyN����Ф���J��E�kd�z��vL��Ok�V�ތ�
?�u��_��ҏ��^�=�����*��fC�ʇ��e�<����Q�@_���%�R,�is��n����O���W��w��;_������d,_���QWcI���,����5�6�q�_��ɳAZ�9�e�Jۙ/˽Y1l��`ه��#=b=p��G�]�dz�_)��|���_��_��*�q�0����M�7�xs����WU��;v����G��7^{e������b�����7߬?g����Af=����Qt��/�+�쩓Å0�'�ngN>���p���õt͝1lX3{x`��a��eòEs��`]�ʲѝ��Ĺ`t�.���C��/�T�0J� 7Z�"�0�m����LC��ұ.�̀T{���Ϛ1�[8?1�J��/�2�ՇaX�����i�tbޛ� �Gݺ�����m�s���x=������{���&6+�}q]U64u��u�U�E��Le)�݊�ay`����E�E����v�4p-�a*����������K�n��ۀ5��d��V�Uby���h�O7��5s-�_I�W"\� �Ev�
I:��t����kf�:]��+�"-n9c2Ws]��r_���Q���^۴���GO���Q��o��i���6ס����n;�HD�y?RB/0G���% �RX��t�Qr-*d���G����y��1V�y��j����2�� "` ���ѝ�Pzb)���'�X�	*���_;��x^�����<p��&,���A�(��k,C���z���P�,�h���k�fB�� <m N	�>Ş��	���޳gOz�G��((FA�aM��.��3�r��2̎U~5����a�9�#�3�֯�����m]?���6�gO���=�n�K�1�ҹX�>sz�D
֦��r����b��J�}/�nX�h�p��M×�z4��=lٰrX�0��mW�P1
�]Hz�#	7�+�Ԯ��,���;|��g��|�������s����ڰm��a��u5���R���Q��Sw�TM5��8�����|��L}1M!���PfNO��0|�<7��������������[C#�:q�V��\�l8w���������aǶ-��a�����h�т���f
|.����U��g�D�n۾�,�O>�\��4�&<�Ѐ��h�(����c���Ĵ����X��c���L����.�=A���v���]�nКU�r\��i�[�������+�+��G=�.۱����NwԌ�t�f�&����A�=@�n1*�I�v¶Y.�>�9�S���eܭ��eC���r�oN,U�@(=g�>F�.]��l`]NرȂ4)�*)K��
HJ��*��1��J���i��5/m�6�,�*e�z%�jg������C�Q��]>�� 
�C�R��QۄԳI7�)N�6á��L>��i�]��78�z�3J ����k��`5�8T圲$?t-��}���5g�Q�1ʵ�R����5��x�ʣ��5V%���9d�-�����(��)�c��������D����q����\hꞺݒ���,���h"�A{^����)�R)3�"6����{�t-��Y}�=�A�deBS�4ۏ�q)��Y�}h˅&oJ���ͯ~N�_�?�|r~8��ݶ-����_~���9�޽�������F�F�T���X�g��a�4s��G�AS���iծ��M�ʭܘ��?e"0���˗,��?��.�;1����)�����:޹u���/1`}t�v�}ߺX�vM�B)#x���e�~�����x�ڐ;7o�����@�����n�Q��,h5Y摇x��(�-���w�Iw۝Ý�6kW�\?>L������1;�V�7�-�6U�_x��ۆ���R	X�n��a�x����G�?��3��qg���db�.�T {��^�Ѡe��p@�E�L��
�=���}��<��n��J�3��9���<3N&q�r(�Ԓ�(��jk�\%�~�����Z{]�r�-�e��-��H�9�3� r�@t���|�sows4��_��{�7���}Nxӆ@����:��\RE�]����S�u���.�I��v2YK�,���⪨���l\ �GCC0
@#"�h�k�u6u�������, H�� =6j���n�0I��`KT(�������������z��v���� ���X� ����i4&��E�o|�v](�� ��F�Әn�Q\��<�*�!�o6�gA�\�Pe���Ċ*���I! �P��s�>�TN���Vj��9A?��3��o�i]w(*�&v[��Oܬ4�o�~�2Fd�Y=�E#ˉ7��ڤ��y&[�������D{����}��;�]T7k���/L�=��sq����lV|HS�|���|�ߟ=H�������([ɇ��C��_c��I�H�2�}�W�	��@�ҁ�̟�;z�H�X�8
��=i?B!���w� ��5y�~�S��L��.m��W�ª���h���ґ��K_|%�x��m�;z=֟�)m��\P{����Yf�O�#����5C��ݏ},����
���(?xڑO|�v�I&��*�o�����J':*7ePsK�˄ߺ�^У�ϐ@��ѣ���1�̹���(��h�Cɒj����u��۹k����~?&"X_z��+ś9	�E�P���Swg��g�ƩOU�28-b�Tb�W˼�XQ�T)ӌ�
�����'gcbVDn뎶��S������^���q����1ai�0ђ�tJ�%�O�&�ލm�;<��6`<]���)���������Nm7��8���}l����H��(�� ����&֧g�U:_�������s�h���ki���i�Lvk�=_kU\쬏�ę���s��2�u/Ǘ��z���������B ��$�x�WDW�F�|�jtx��F����LZJ�~���j�_��������w��Ҝ�T��ۦ2�<<�=V+db��ߢu (ۇ^���f����t�p.y#	y�(���7@��U:�~g3����p!=4u�X�/�;��Ơ�3���l�
�h|<+�q�6�f0�� xxϺJ���y<��6B[����y ��tU}�G�!}�ɫZy�7�M���y���w�wݩvO60ρm7me�/�VI6�ǂ��]
\� 2���W��_���a�I!�	Z���]��z�(#�<�Ze�a؄���\RVY�|�G��L�;�|��5h�gϝ�
�l�r��U���7��0��eZ&����K��Â��O�O���T��14t z{��,�W/k�q	�.O�������kDI�ʺg��*D-�H��aQ���`<T��{0�kq����8��R�hQ��?�Sw��.(�Jp߁��cאv-�|����Į={��n�O��j�6zwEGw{�-nħ瘄u'���Fخ�{�!��0�������3��L��
�Sٮ�dzkxu�v%�&tF�շ�äϋ�D�����dƸ.���R����F'�P���8X�0oln!�<�t/��?v����g��Z�*w��.��������lP#A ?�߼�P��з�=�#�̳ �g���������Z��kϣ=��<+��p@ ������ G*
����Ic��4JU�~��f�%^}G}�s����7�E�!_X
��A�|d���+}˵�+�H#���q��y�o�'5��b"��i�h���ՋT̪�j�oKm��^
�f�f,?�L(�M���C�������5X��`�Z.9��R/�# b���� ��7epBC.�� ���)ab�vn���������C���ߠO��3 !�W�J���(#|e�յ�䗲��=�fq���-�h׉�g@j��o�g�+�R�l��ߴ;x��@ #l���K��W������җ������ve�+�Z�@g埶���M����	7R*���s$a�[�!^�$_��ˮo���02�WOpP?���|�\���RM�G8�P��`���q��c񕯼)�7���S�⑃t3�q���^ӟ���LeOsV�= +�>���n9�7&��H"u�k�e!��ɠ#�oF�w~�/s��R<�����jꏚ�V/��jo;v���6�_����\�;��舊��%�.�UI4�a��3Q�m�Tx|݌"��bX2�a	��ĕ�*��	��|	��z�0b�dr�͆�eKܿ�cuz=I͘����y!��:�6���Ko5yCD�/�1�l_y��x��/�~[f*>�\�4AfH�U,E@��x��3���o����^�g�LJ��9��&0;պ�3�ę4J�Ȁ%@@8 �̶ft�=,�Đ\��U=[^��V]���.8_�p�w��$�L��N�jmc�6��{��hЖ�&^��kj1A�sZy�F�<|.C����ǀ�k~r�K�-���򥌃��k��t����.��@�!���t�`��^�� Fz ���V� n	�޲S ��x.|Knt>��C�<HIS����4��Lq$�R�%&�
�A�|�?�����}ށ��C��{�^v5��bY練���_�	��p�v�f�(��͛����I����s[�*wֻlS������\�zМw�3G��X9�Q��0�cbm?��������m �z���1�&?��yS��#���d�1�Q�6j��/K�O^��O���p�r����9�P�R}m��@��H� �H�Ι+�KgϞ}^���W�(�\��d?~2�x}��^/GϦD���{��f���!����w�~a؂����e(&��ǯ����~V�c���R�g��娓��c�2#	20��cJ`�,����kM���?�ti��WV��-�$�Xʘ��LĢ�������`_���s4L�� o����X���h%z7Gd�m�#��������{v������T�?w�����3c���G�ƥk7�c'�M��3����3���_��ŀ��S�<��M^@4
�=:bX��Nm&�--a*�GB�I��l]1�!k������B�� �|�3{���ri,)Mz�o��r�ⰖF'/3���`�fK&��[(��s/�t7�]:׉�F)�#� k���S��?W�E@�g�;��aF����|!X���*s������n}*��֙o�e�x��-��&x�y.�>�X^ ��Qi��O�f
�-}p �|��D h`�-��gh���Ψq�60��c����M�t@A8�Ec;��xxz��y��K\jkb
�����@���}�0�h_
�����г��i �]J���R.�ǻ���y��/�Tf��'�P	� $ k�U|�;���GyQ�2=��t��f�J������
��AY�_y����W_�_a~�.f�	�(gҹ(�x�<"D�4{�A�a���.�8��g��}D|�Yfޫh�Z@�cc�G��0�V��m,���;��v[H,3���§\
�%�{z=Գ��N�~3.�-�������`R+�}�k������Z�O%%���t+Q�������g���;�ںD�o`h�9����������8�^�ή�]����uaX��FzVW�b��بTC�U�e0����Mà�1!L�Yc��!���z�>f�2�	]���g�Υ�}W�"EKs�U?��3�7^���F�_�2f&��^Ȧ�24���� ��t�f����b�=x8�:�����8s�b�����o~-~��;����Wd��H�\S��H�P�q��ӥ�*[!��o�`e��� s"�M��ǽ�|��	f䠱���	�,�J�!P����
 K�08Ze�M����v���-iL��-���/��H@H��Y��Ge0�km] 'ӕ���uiz� �i$�0��A��;Ӆ���Sq�79!��f���T9t�==ĵ�	O~|������C}��ͯݖ ;�}|���?�|�9��T�賡_��@�8��^ �����Қ�e�_�2h��:GR%�ܣ���o�f.^eR�ܗ���/g#�@�[��q�p�n��y o��/&�hU
K��Y鑦����ɳZ�-$i��M���Ƥ�Y���A��i�Z߃��c���Z�ʂuE�L�b��i�zhU����2�jhl��YP�Qܫ���G�_����/=oPg\����N4V�I3�q�,*�,� �
��mD}�J�i�1 L������P--UY�Rv8�͏��?}&%8⭷?����[qY`��g�_6Hb�(�}yL��wך���c��60bӥEa�1a��Yb�V	��v��y����L1q��M����� m�����X.����
���OLĝ�[q����;�b�ӌo��5=�w�N ��A�����:"I�b]&P1S��3�"��]�24U �R��v�u�>�N��Him ��h�FM�m!էƉ[�ʌ��ut�����5T�>�2z���7k�/���?�ƭ[�,�̬1��FZ�q	�b���� /<�t=��۵s@�[��X�!S��=�ߗa@����ɘ�=8з-�;0���M�;��p�@C �º�ꝕk!�(Vk��a+݇���."�kj��`|��{��5�4z��W��j�u��1��I��Lg�6a�Bν�
]>��73��NG:}(]���~��z�g���h72L��7|�����iF����_n�F�K���@���C�D4�Y��rO6������ߦ�C[4��G�OM��Y�@��"(q� ����P�X8������_gx퐸/Ʒ[#�w���9Z�� �� L���a�}���{��p�������Ѐm>˧����yV(y�7�����U��#ޡ?�<3���rR(�E�]n��Bm̛�PXDt�3J��,���(9|�V��;c�J��#/�k_|Y`�dl�]o��u�Շ���O
��( ��>]�޵r�#��w�74�Oвd^J�D
�`C�������C��,�����7��y�>@h��X�bD�;<|[�Ԙq~��z��&���1=�'�(:���<3�����/\�X]��>���?��r{(�^`����;�j�=��g�^�9�����E ���4��F��vf�<@�hmI�|�] ����jؘ[���"!�7�Bw@�	\�0�`w�H
-�$x�她&&��v������@b*s����UF��)��\���o|�w���_�`4.\�O?�\�޻׫c�9��vL�V���^~�H|�I�yd�Β����y���e:H��(}� ���p��8�r�o��D/�$�{g]��`g�W�Z��.CS~� ��$d���=�G��Ui��Be�#�[�(�Xi��A��d�)|��`͒YXj���9C�r�a��9�fDg)��t�$'�#I3`�x�f�s�p�9����?0��Ͼd�tA�E����r� ~�Y�#k�Q&�}	�pT	��E���Aqϝo��K�ݎ���G\<�6؇� ���Y��<��Fhhܧ��I�����A�~���6�wy��p�?s|޽�; ��M��^�-Վ�j�Kg�X ��Y��w)��h�����t�0{-��z`��ˢ2� @_�)k�0�t�,�(Ї��Up[�r� F~0�rQ
++���~��W�o����4�U��M�� �g��QV����*N"yƢ��A8��Ptk ^"��;�)���J� ~_�Z�u��Xvt�/x)�|x�1�К���v�Ņ���P� s��J���ܭ���~A�Ya��tzd�Nq���bT}��?� ^	nn&禣r}UZ�4�E�;]�UbZF��Kz�A�lR�5L�Y^�
�p��G��ާ������{��Y ��(*�HSҕ�6*Xt��M�A���_ �ށ�ԇ5I4��b#��I��b�$%*�Ch4(&�0ĊsW�@4�v�3Ͻ�%�/\��/�sG�xTcx�Y
�Ǥ"�9:�Z���p�뭛��ԉcq�����Ը�#�M�ܜ�V71��V�i�LI�}+�]�Ο��z*�~z��ӧN�'����gϺB���^�A������Њ��{ʺ��<%~�+0���q����x�]x�N�O?9�Μ���/:OS��Mȳ�����@.��A47��y���x��=���KGc��!YS9z\��2�&M#Ȑ� l?��+�n��k��($�A?�[4P�y
mB�q�  �������p�}���^��,X)$�Z��@��"H'�.�7�Z�� 0 �Eg4\��(]A��ȫ�<2�i�L�*�: 4�$~�����@�,#gǘ�a�(�o�?�yG�6��_^v���34U\5%�گ� 3�%��\����,}ګ�d
��VOw�-D��\qvآ���ٿ�xDn�hߊ�ޥ���4���|�l�	 cu���s�wh��{�M&����P��_�O���i?��4T�� /��H��M�QG|���S�%��+��{5׶v}�0����9<wFG���ͨ�KA����γ�ޔ���[ᝲ�;;��nmV�r-�a�8gf�2��a�,"��ζ��?xݦ.�������}�����_l��R�]2����$9�LV��h��o*�Sf�'D�7���[�&*Z��Kq���8}���5�ze��Xb �Xe�B�v�@A��y��~Bő>g @�@	wRs�'-xr|,:T�W^z!~��7�)_�S{v�k���Mݯ_�,F��`75�GcsG4�tƕ���o����_�*��?�W������G������l���^�as������w��mM1v�4��x�����h���ۢZ!��hج���M����Q	��\�F���� K@��hllD�Pe��zb�����Hw�3:�.uR�0���H��E:vO�{�`�|��=�l|���35yx�1�t�)<����]�����/�z�k}�ߌ���w��ͱ�����x����(�S�*�m�$��%�s�Cy��M��2����w�=ɏ��S�z>DYp�U9 W@��] �կ�]j0��<�N�P��<��]�ƀ�G�� f3�F\�v�� B��h쯾��wp��s�+�,q�W�,ꋎ��~��t0�p`��C	F��&���p��iB�Ё߸��ν)4�2�|�( ������5�EU�9ʻ���~�	aT��yLi@?����_|��	�����PJ�)��
|O����s�}_�g�2o�4Z�~�Їw�c�;��GF�T����=q���8�  ���/]�bw�W�x=���o��'S�l�"���a�B�ץu;�S�O�j���	1��t}y��:u��_�kkɖ��=\�h�$�a͡Ç�~)�0�^���^Ty'���D�.�Y�d���*n"�\X� c��_>*~S=��ʶ`!i���?�9�A�H�:q�W�ߪ�o�F�����\�����Q����(�@��#�Ďގس�/��ޡ�@ػ+v��L�C����=���C;��l���ث8����;���w�ꑘ6��5*bHW�#�H���h��z����OS�����,4>�PaaQ���k�N/��<"	�F�r�hhS������S��&S��<�q���p�R���s/�\��z���{0.���ՀϜD�?~�n�>���^ы�M,o1'MyV�1�y�π/ ¤eR����+�e\�tn4Т����P2���+��3>}��.�=�����{�f_�L:�q�0��F��~��;�;���n��*3��*XjP��Kt�U�������\����.�
�I�i�0X�	3v͆���]�dY'rpd���-�������[hs4�R�@ý{��+/�+�WJ�[n�G,~	�.�IM8]5�	� dq ĩ{w|�q�ŷhS�]@�ƈ�p� 7m �!OPR�4T4d�K����Kڠ9���yh$�2�O��z�4�"�2��(5�dŠ��	PG�wP{���_Z������C�QF��Qڸ$H��`�xs����q� �}|�X�O��=�ޗݑ�.?�7�m�����%.h��M�ȵ��-Ęi���C�ԓ��� QO�R�i�w݊6�Mt��툶��|�g��)!��=�E��� ?���A������Y����
v�c� ;����}��gm2��\y��i�@Iխ�uѢssC�����D�fi��U����R��/Y;��[��Bq��S���Ʌ��w����?�<�1���ڪG��&�[DJ}�ۆ��	\<jb2�1�] �3���>g��'z"��>6a�{z���5�- ���}���h[�7����L�υ�kH��c�Z3=������{q������'u���`;C6?y�L�=w!N��Ԯ����xIZݾ��%��{�d�Ek��m�GN�,�v�,[�`�ʴbs���嘞`��q3���m�� B�g4:l��Kہ�=�.�a����,;�9�e������{��������k��
X��מ(&�`0ٕ�c�'���b%0��NMU��5b\0�Fnܼep���g�uC����/�W��Z_S� �Ͳ����hx�*���p�T<6ϕ_ ���� u'�=���=�(�@�ɉ��N>J�!�r��E��� FY�� 	x�2�a����s�=���]]6��%� -��'�' 8��(����Й ���"(�'����] �b�-ф{��lU�>�l"���T� &,U����>Z-��4�f��n����&ms��=4����8�������%���#�e����
 @3o!��tx�v���|P���?!�}�JVC9O�����>+5d��e�Y`��
R��Arɴ|�s4| ��g�śmR�zd5�K����<o߉�R|�����^x�F�u�y��1Jp��{�.}[�*U&��� ȱ��6�x��T������s�0v2~���~� `]�Z�+2�g֗�a�M���D,Ό�܄̴����t����z6�O�|Y��չ�X[��-J�	?�Ҹ�*ј�AAS��L�9���A��ꩢ=T��a����I��ߖ��y��w��M����}��/ގ��^���{�ӿ���O����/ߎ��;q��iE��a9�f�w��X��nՏ��f�hWh�9*�jHt���r�̒������]�p.�{����/~'O�K������+5��F1.~S:ӹ�QN���b�<�z�T�c���K���>�s_y�73�K�w��� �ߵc���##����cq��Gq��E	�I��;�Ѐ)5���|{ؘ��e'% �M��nN�Fb3ZR��&�v{�|��͙�>�����{[��Z���ӝ�A# /�퓿�ym�- ��D	7�|�p�۲qI��. �ڵ�o�E���¹t������k��qc�I�FA���Ё|X�����<
I�Б�k��
�ֲ�"h#��E����.w��XP 0ZX)( �G�r
h�#�#Y.�Ÿx�c�',�L��rN��n�,>|�_x�v�m?t�P��a\;�@p����ȨR��x��إw��9Y��Q('ˮ �!#:B@@� ә8=Im�a�̖�A;U��^išT��~���/��x�9�:4�~�l[�2�}�Ƀ��V�pM���ȣ	�vj��s��kL<�AO�O���SQˬ�u��OՖ*u"v}�ـ���/ߡ;�VqMv��#�����Gh5=]��Z�bj�5$'�t<pƔ��X�Ƚˀ�
 ��R�/��BM��{�L����H���u�"�l5B�l��r��<��<�c�� ��^�D�M� ^�Y���A|@���s���+�~�L�n�oi�f��߬i��7�N�W_���7�,��}kٝ���j w*��!t�6 ��T�U�R�n�  �Q1s=�P�:ٿ���Ξ9�|a">�%4�ҩ�)��0�P�  -�IyS؉I����x�1���)����j����-+>���!C����A>�������,��'OH@]��裉��]J���HS�.m����h8���8���c	�50��M�Q�Nެ��S��M�͓��yʲ�}�յ.��nnб�q���#�pװ:'��AA����8� �֧�� �`h-&9� ీP�P��9b�*�~]��.0�:�7��8��Ra+ЀCZ�]ֿ'�� @�� �d-_7���ɌB@� P��ӆ�P���q����C��ٔ8�x�x����d�LڦG��q���b��'�x"xH�>[9�8 l�!�m�D�6�>#y��E(��8Їﰒ�z�l���b^V|К ݱRHc?�|:��(���}�����p���W�K[N�?�a�&aA�K�V��u�c�9r��b��E{��S���^�'i����{qs�n�-�(OX�?�	�Z(n\=��w����o�<5E=81�M�\6����F��*��b"�}t,�������G���������R�L�Cxk$�Ga9 ��7J^V�duIZw�*`n~I��0F�ƣFZ�w��s�F�ٍA��4^]귁�`�t&��D�!�����:� ���M�߿7�~��x��W������3�<G��/��E�kq�ŗ��_�#G_��_8O?�|<�D��օ��qA�?�W'P"�`z�=�ft�2Ҧ��>֋Ꮨ����n 4ď>�Ȯ&��"diȔ����E!%d��U�p��,5?hLd���:C{w�
�tS]4��X���̧��ܓ�DP�pZ�9Uۯ
���3gb�����4\�́�A��Ff	X���ݸa>���;��xf�Y\̃(w�*5,�,���"��#����8�̐7�^�t��)C|��^"���h�칋Ϝ�d��c��]�A}pxy��5��`�<Ѝl��E�&8��t�d��΀,���S�ċ˂t�oʮ���|���:�L[�����ƪ�� (�>��$����3��;���q����C�`�X��5�<��6�@���g��vi�M|�䉲cQ0  k�}�!�@�E��
���_8o�C�y���:,���"/y�����51I�x���}{��e��za� ��[�M��v�-�`�TP2�~�����o �-��>~�����!5�`�����w�:��۸��ÜUo�����\�;42b����Xpm���x9
�'��=QH�O��5VFZ�[�Y�����Q����ƿs�K̑���b2�����&��i��� nLf\ʡ�!��['v~9ňBUM�g����Y��4D����ϙ���J<�66�!3o�o�'>A�Q[�*a@=��]3+ SΪ�`b��`���ƺ�0�����0�8�Ͳ}#c��ah�;sٔ�!T�į�!@��EҖaS�7Ѭ/]�'N�#?0��ud8$t�w�eX]F�T	�0:��&��&�=,�2�#xe>�8�~!~V�C�>�L�t%��@H��������B�1����m4N,�/�ұh���W���=���:�I��@ʺC�e�2O�
������o��|J�O�H�Ƭ� )4��ǥ	���㧱� �ӰF_ąUF~R�"@ߤ�
�B9���p��zr��gY.\���ԧ�yXs�����+i�9��u���~Q6��BZ��3�&�� |�f.��w=n�w����^���S���rŻK��py D��w mh��j�h�0�hd8nɺ�7�0��#�+�L:��腢��U��21$e��KC�N*�@��zB�&��%�#��24�+����m-Vv�k��*�T^]Q�0�El-EX�2�7�o���)P^�ߕ|��R�h�A���E�͞������.�����ǵ�#~00�zA�i�<��t�����W�5~�v���']h|S
�!�#������\��'�r�����/������M۔$)�[%5(N�=ؐ@����P��?)�����g[4�m�� ��c�I�����	<"j�����k]��ݸ�D,][#V� �1]o�o޼ׯ]�˗.�ŋ��ڵk2)G�x�mi��d�f�]�|5.^���\�y~#Ν��M؀���%�����1bA\�a-�3|��j�-�2W��?V�X��,S�ˡ��.,��3�ⲡP67T1!�0`B���J�@7hķ��x�f-L$��`% ��Y���|�{^g]��)���T㤣��y�g��m�MB��<{��,��7����>�y`B��Ty�j�;y���yl��vPv�[*q���K@d{D3���9Y�������1�A��8��U�<g�V��A�u!ک�4x׏��ڠ�3t�����H��������� ��,��ڂEu���������g�3~_�r�'�Y!�]��3ѮH�gX�}hX\Cg���]��x �0b@���6j�B���.�,KK���={��a!<x����>4Gp`��*�ӞvB��4h�h>�~F�a�e��:A�Ț5�8��ޥ������3�"�fH�2�:1�	78���C��wvtʢk͙�V��}��-�^<��uЬ|	����ў|0��!�%�a4~��4���Fy=�~��;VjX>˜�u� ��z��x��*	 CĘ��GW�T/����Uw��u�و�e��P)xމ���,��b �_Ɔ�I���@�33��EU��|�7���E�Pr���^q?���.�4�(�~ ��0UZ�%�?���x����U���cq��Ÿp�J�9sA���x����wދw�y?������ǒ�'�����X�֖6QLPF������nWied����3lT���=�XxF'�?�P8�[0l�hht��φ(��`Z7h��!uH��]�s6 }B
73��Ns�lz�F���j�G����e������䨪L�Ꚅ�����Rf�86�`�-+��;�W�E���>����]
Q�~�=�ә�#���e�����
�<���@����L8�)����#�� ���i� (Hϝ��'��� ����G������􉏃��U���9�K������� Q���I���[�c�
�V�����C�&/�����t� ^� +�,7iCO���/}a;����]S6����`M;�6�UZC���	� ���B���ʻ��`��D6⺴��.�C�AI p��ي�7%��	G�^��W��'y���7i/�?��⫰�)�oX��39*ʽL�����B�2õ�2;,wR�uE��.��m`u�zr���q�$*�=U��ӯQ��m��������0�Z�=4I*��52� ~��f�b��`l4���Q�$2�7%�`֯KI1yC1�WMUY���o�\诤2%��G�=+�nE%}��0o(H"E$��eq����#	-�Z2���$cCs�7wDmc�Cc����+T�U�a��d5R���j��3˓IO5j�T=U�$��TÚ�� M���d	<������x��
�L�f�V�*��ǹ��Õp��҄�}{'@&C�)�h��@�)�q����3�	,�����7�o��%�9�Wx4L�-}�0�4�k���\xG[�������.�o(a�
U�֮�MrMql��~�'e��w���Hh4�������D��O��M<Ӻ�7 ��-�U]q-��=@���&ь~������ሲ�T����rd�$+3.�~Yr1�7�OH����|�fi�91�޾��	� ��Ǻ+����#�M�G�	��[@0f�}��B)[�_����7��Ț�('�!�"��N;�]���>�I��e��{�yw�J)�U>�X�U�X�C�CwH�o��S��8�����4��?ިv�8Ua)8p���+˸�h����= ,���*>��L���5v�S���@}m]��Rװ2�*��� ���֢O#B!q��v���39L K4SV�h�������~(B��x��a),f�3����|��ɺTw�x� �-J�(Z��g{��\H��g�i�$��e�3j�aK]��.%�=]2�w�� =�}�����};vEK�vtEs[�78awy*�ZB �`^`<_�� ,���I����\A�Lc|_���u1��!�H��~i^�@HY4RV��1����.�d�4��U����\u�Q��U)_�
��$Ě{����Wϻ�^��[e���F�L�	��f�e�(��KM�U j�
fJҤ�`*1"�ifiV5�%�8��+z6=;'{��0^z�����������,}�0��(� ��Ў�������}�2͟I>ҬdQ5�seU�hx�� �UY�k�Z�Q��� �R�( Lnf���;�u���2�ŭ��I�f�+�F��y��K3���e�����Z;�� ��qJ�̨xTL��	�N�jɮhG �	�����#��U^q�	F�4��^B���XP�5?���xJ��&�;���R ��v��V�Ɔk��akJ�ڳ2��  ��z�N� (k�J�>%���0GУ8xBўr�~̱,lcZ�Y�?�Ƕut( �-v����/�U^����V����t}���=��#Z���X1�?�v�@^F�5���9 �*U@�I! ����c�㠔����(B6iW�db� Z�����YKC���4kT�ц:�M4�F�%Z17���W�bt�AܺuGϕ�~���	LU��SIL�>;k#�"�+tƻ�HmO ��	��	̺�Ŋޛ�����%����U����F����Bx#�ᘟY��#�q�ν��u	KX�rE�������:��F����3���xN¾��,DSc��t���;��ݕ;�>=�|f:�ݏŹ}Mu��^|V�rUZ���㊈�VH�j�1��F5f�vv2�]ɢ\����ho�uu�[\�_��9G�� i�S��%L�e��2@���Ր+D��CЕ���)+Pܨ�4tFۧ�`CL]!��c<�5`�����sf+�ui,*�#��*鼢��U�+JoU�>ҽ�Z 0��HC���!m'�Kv��Yiص�4)&*��Y��̈4�-A�Y��GsS%�(�� 	����f�N]��Sz���l�s�3h��i�2d�+uzw�����f��
��3�ͼ\�
a��a׃�A�+ MA5���
��"zo�"��6�2@W��_�M�O_AeϳbV�9)z�?��X.ʗ�aj�X>������r 3���S���E	e:�M#	�8�
�=�EW>e� � �������20v��p`M��y6�,�(E����T̕�-��at��X閂�֧��8�H r�_g~�m�KpO����eg&g
@��^ğ�(��2X��~��gH�˚h�Ъ�����+���O�Q�Pj�5���Q����&� �Bv�>�b��Ҫ�hQ�k<p��Knܸ�gyZ$4�_�NXF�s./m,P�@�_[׵�
ײ��M�X��zL�X�$!���Ż�����>��(�H�%��M;Dy�������|ak<,�@�`�&��ʏJ��?�l�<I�02���U1z�a�-���k���"`"J�[�⣥T�5�2��m%�d%��)A�!B֟�D�I	Ӂ��L�w����CŹT	�����FP^2
�%���\� �-1A����ξG9�����"����1�>�iD(������gI'Q�N:hr1��� �Hp9���R#�kW.{�
����YA��k�V��"%�斈f긲�;])z���μ���<�ė�&��(��{�q��i5�32�<t���>�[Z,.�#+����ШZ4�;���#�4���H�m@j���E/��W�3w[�j?���|���ߤA��k��Y��a���s�_.�Ӵ��3;��.=�� |���8�]��O��������$>րa  �ݱ�CH���h��65P�٫���U�J�hpm<W`~#�H�����<@ï�wLOj�O�+a�-���Q���:�C�G�m�:aS�z��:��z�ϋ6�Y|�Nl��v�CI�������F�0��]��`����2��\g�.�cB# �(ad���(,�:EUa�"�ARҰ0HT*.�+��-��j�t�Z�f�$Y������]�+�gv���YY)ZJ�S�*��x�/�t�5��[��2�x���ĵ�{�JgC��]Ҿ��S��d3�� �ã��e]��v�F#"����7;�	��}���8��1����XizY}y7�z��m�"r�?/{���a(@߄ )S0��Xub�9�?�n�Dub<��A�8�ag�e�M9 d�u(��5M��(�%h�s��ٷ��,�}���6;;�S����09���;wy]��2%R9n(����5�-hԜ�v��`Ν�OO��׮zM1Z@����y�7e�� �qҥ�sv(���o�P|n��]?`N7\�H�g9gf�޺Ų7����ؽ`�2꿏}��q6K:���\�HLUk�?�o�xM�������-�'G��l{����=�vvE?+�^Q�ȓ}�E
t���*Mz:3���g`��=��8����94��,@U����Вk�,�&��/�¼I��UEG�>2���5(~@�MZ[;��HVa����#�'h#�߮��n�J!��2��V�Y��Է"��3�3g�KJ��v�w��#���k<5�r�ճh].̦?,������;~*�V����kLE��L:�;��U�����Hps d�R�X ����]A*Lܓ��ɧ����7�Z�V���:)+"W,���3W�-���֊��c�7��V��AɱP�3^~q��Jl8�4j+�������u��l��W�$>����#1��a,J�T�� �.�p$�I[�n�� �4s9u������- �p�1��tR�' �֝��1�u\:C���5@�?Ef��JN` xX�}z�E��<i�����8Z�AE��o�� h ��J�$�b<�#�Z��2����Q**�|���ˇKʑi�����3L~qC(�v0��9C@�5P�|���eR�(k�g��Y��-���8g��*�,��":�D�w����q����51�Nc�vhx�h�@�i:�W��Ժ�i���^���|BKΔmY �&r3����ԥ����ݷ�k���zz��e�;zǦ�2���"�?�Z���F~(:m���yV>���,�#�Z'��w�3��}��	�R~ӊxw	 /��3���G���YW��u�$���J�����@\�$��:��f;�N�E0 d�{�ro�K] #4nh���Qn�'��}����ֺ<��K��~*H��\vC?w.]@���	��͟
�e�.*���6L��I��:���~y�w|�+�����:�#J~*5dnE�������mIY�n�%0<��V����ʾ�Ds� �:ݧo���+sI@�F�(i��U1���W�~�	O�$X���i�F��Z���P�K�iU�)Q�^�C.%)j�'��bv=�3M�
����)�s#X2y`G��uKӗլ�s߀xQ��r�V\�)�jD���`_sq��F*E+�W(�����n�yŽ��"�t�a�`�(p�������#0Eq�]\�.�̦�|9C5׻���������০ƃ��WfޫU�����(pf��3L%��l���ʕ�B�T3A�2�ϖ�Қ]�dsA ؂.�s�O�f��J��Io*r��N��GB�p�>~H1���I�Ȝw%n�W~��'������9�%XZXL��j��^{�����ySt[�V�6��$M�hd�Ng�z�٬���:Ia�o�t���x�� I��4��
�=�2����Y��gx!�4��ߙI"tN�?�d'>���'��L���}�&��e�)Z 7gs !��^�<���h�z��k�آs���yؚBnC���z�3����~�_wJ��}i���x����P�ӑu�Y�}d䮬��f��q���zz�3f�s:ˉ�@=���z�Dh�h��%�Z0<��i��ϘDg�@�]'h�L����c�z�����D&�<Z=@o�Q�I[;�Dۣ��+���wvw*t8p��3���4Xp�QJL�bl:��I��`�*��5�n�\�;͔a���.�of+5��Z%(�}�9�9@�����}k5�zP��.����������w(�Ш�o�ɹ��������y���4�/�.����R ����ɇ��1Y�V��d���/�7K���<|p_�<�t��JP�J�oko������\���|����l�㟜�[w�bEy�kj�j	�G�&ؤ�\�x����'����;�S�O�;&����q�,�ơ�0_�}G�SA ���#�?) ����~Dd���!&'t1%�vы��� a�� 늳�;>R�^*��Lp~vVRq�#�2S3ʠ��ؤ&�P���{!'��0-k
4w��{�Sc ������T@�y\�@�Ǝ �t��_=
�+�~�8u �R�i����g]��tO>�Ly��U�S���L� �ďo�bX��)�5:�ʎ6�%���H�p)��f�6��P.L��^f���O���>����c�UvLx*=4Hm����8��w�Ug�xf벸�^و�<���u�n��Z=�-�����QJ��sG ��=�1�W0(;!�?�=��L��M��=S���N��|�t�&��X���ǃa��DfUV	��%�	���,3e�9>����*���Ĕì4Mw����Q��f�u�upt�v�o4G�cY�-�*��<���t0�:;KU��%H�g����:cmp�ݩ�>�t����7	:��X� g�� `�U5��|�ss#3���e�&R]XcTڞ'�����V�����uè"�s_�w�=��!����RcX��`$�Z��G�бK[Y��J�
u���`��\:Mw<S�e��B�0g5�y���\�"�%�}\����!���90�;v퐀�r�tR�v{g����M�:���d�M���ꛣ���J�C��L�"V>�z/6$̛bߞ]q���Pr��
8Pb�	�+MI��)��)F���@?�OX�hnnU`H�����L;v<��������1�"�&�޸D�MQEJ#p�cN�%1%�\a4B5j$}!$����"��ꘜY��4�LI�	���V6)E�>�<BHKB������� ����v#�W�|#7tbX��t��LV=#M���R~�c�T�|��Ǣ��ǽ�&�Q���9����7?/�(-�cH�G��L�<�qT�rde �L~+���]��&�h4\��[��G)��8r���r����"� 5
1����I�� ��z�A����D������ᙀ7���Lc=p�عk�r�{���H�+J��:$E�$N׫�Ĩ-I�" �E]C���OޕׂVz��*}�v�����_��g���!��DS��d)�n�ƈk�ۂ�a�efc7�T��kFp��wH�H�%(����m�5�أB�-�M �,@@��uy^X�3=�7��;! �Ah�ε+n���q�zw;��Y�p�xCP�x��%�
8+����3�93�hYH�w��yK)G@��h/�e���S� �N�����N�A��.��f�Ю�i�E+�kD/���  ya譒�v��[��j��%������V��sX (?����^���,�Č��%��rq��W7m�}:d1Gc����:�^X}�d�QӪ:\����{��+7��꺄�@e�QD�@�aŢu� R&�?6Co�����%JG�痾�:���Vy��h�t�2��EIC ×�'^,���?������ύ51ˋG��Ï�kW.J�M�DE�h�5���$�g�6�S��(�/�d����'+�d2?��.�'��%�;bm�:VD|p�9C�r[A PŔ0��V' ��%d0�����nЀr�g4&��R ���RI�y�ʳf������BTn,GwK��|;vt�ʼ��������i���3g� J����2"�ܗ�9)IM��ͤ��t�D�Lc%q�4n�r�i�k��nXkWY(cY.hE��=~��ŗҸ��->MFn`�WZ�A�!��2����K-�s�8Ѧz���;������_�'?9�F�ƛ�G^|%�
�����,��{ᅕG��ʛ�Y@U�[���W�z�w˒Ј��|Cg'�&�q�M���ߍ��|B�tܾ}Kܔ�L?tB�� �~_&J<И3V��� �!r�R?hn�2�W�\��lfj���/�_l�U�/m���D]Q���Hb%B|km_�$6�)�^��2@�\><�]� +�Lʙ�:x^���u�Eޣ|�v��t� :��k/� �+�!y.��4Q8�͂Z@�|(r�:�?�[���uxdY+N�-a}��λ,�E i� �n����O;{wƗ��R|���=�JW4ﳞ�,0��gO��R��W[~�S�x렶�Z�BVOs��m0_���t �nb�KU�J�ӷׯߊ���M����1�,��Ȝ)>�B,�
����$�`o�Gk�ʋ�d�j���o��J|�_��z�G�����)3D@�f�4��?��V  �Z۰�Z��i�OН�⅑������/����wۺu���Yi�bN�^x�(���
2@�T���i�b�0Og��IBWJK�52r!N�������~ʾ11�>Pf�y�"t&^k�R�q���#S�v�E�V��|��L�'��������F�p������ݭ�G?����+V���ђ�A�� XK�h!(]G*���%K���=�S�!Z�x�t=*FYa���!���E�F=ti�B�d�>�!�Dʤ���4�s��@��g��gbJ���y�y)h3&h�Х�{0�>�T���b���?��'N������F<���~��8y��M�RM��4�4������PY�/�����ߣ��}+�l?�-: �hq,�����?��J3/S�\c��t�ӑ]���>�A0sN�\q����{�q}������{q�x���^��1�2�mH�x8����B�g�S^�7��ׂ���:�9��C��n<~��8|`������[ŷ�!�̼Q�#��zZ�6��M/ ~�m�w�F!�O�o�o���}�F�(;�ca��I�L��X��:�g�V0ۓ2�4)<��C�����W�l)UU�6έX�+��;�/����ߋ����}����G�dTgɃX�[�3SM��UK�����|� ���s_TI1jh��
YdW��kߙ��؉8w�VtEmc��0�	}Lr��3v1�ɚ*v��{��Ʒ��F4KwU��g�-M�`ŭC�a�`T#�(5i_#,H�s�.ǅ���������&��.\l>+@���  �JE�m�|f*��J1�)t��ϩ�7��u�S�qⓋ�щ�m�� ���Z\Ɏ5��[���bu�9`�<�<�@��[�R^o�W2=e5#�X���+W�;�x�?*�528�T_N����եYeo9v�w�w�k1�Ӫ������?���E5VLu�W�dj�5�l@��=1>)�*F����`��Y�
�ōB�������1��,�"�  ���c�u�E�S�*����7S	鱢`_�+��bp`��顴��3��e-v#3�������O-�_�?�o�<����%����~�V;~�.�z� ��O�s݈h�ɦ��<����) ]W�s�|W��Y����>/�M����v�����9�+�=�����<&�����Aqp/iU�K߽��+��S_��̖�S�	� $%!��l�-8��}�EH�w��G�y������>��l�<�uTĕJ�ա{N������Fe�׬��~
�x�j��O=�7 xQ��i^�BH7��OYj�!���@�~�` Ę�(�`�[�q�R�$��e)V�)ڣ0��R W�<_����ll{���q����٢�Z���#Ҋ�7�[@�0�W�%nE Zam,+ʟ`�����#j�ţ�JpyR���e�ݐ�e�ӳc�;vq��]�K���X�L\ݐ�(SRy����7��z|�ͣ�(X㑬
�mH/��b�GV���~͡V���q?��O=�M�'��s��+��hF��� �@��Ph�h	����W���/FLű���by]&Ik��V/3���AQ�B��J�\�B%��4ɪ
�F��Y�����(�F/��x2�/g���ӈI�<��	x^/�oU&��E������%�af2��W�]썆:6fɥ�eG�Gs�aRK#�4uY}��}����,O��0}� ���²d�S~����\D��\ҥF�� hi�FC�L�*G�tww�3�e��O`��K���0
���#�z��8��yoT���ܵ;����<���������ҕk��7��:7��Z�/�a�z  hIDAT_��θ���-�����S�W����QB��P��(�Y���Ya�1iRԱ���WZ|y�K�}����+=/�(A��}�{���ʲ�������w�w����g��?����:���g��%����9��Źyln�b!���)���9����qn��ʖe�ӳ��q[�,�p�y(��K:�6ԏ�w:�;3��G�-y!�u����(�:���U��|�Qā�N��S���Y_�6��.�}����g��'�8;�����x�, �Yꠜ|�@a�.4,a��������1|�A\�q7Ξ�7o��@�Ǫ�`�ki�g{w����H�ЮV��RQ(ח�{�w��Z|���B�**�k�������8������Kw���CT��'�A����=C�=V����3�h 5�����]	���/��� �C��_�Y��������8q�b�<���ء��+�������!�< }��\g���y���g��	�����B cw�*�5��Y�-2��x���L��,�@oG�W���4���y�b\�pV����}t�f�=�h�Y�>yc��?|8�M+x�I�t��i]V^y�_����#����=��j�_#�߀:%o�_-��f6�nv���w!H{S�� ����v�oǽ�������o��~��q��H��~�8&�g7��;(}���:�~�7�)��Y:�PQĬ�<xJe���.7�U���|�5����O<h�Y%����T��%?�k��}�q��x�u���Ȣ5>>d?W �ԉ������|���
I�l'���W|S�W��b�K��B<�.N������f��L����ٱX(0	E]e1�#Km!�@<�&]ʉ+�:gd���w�z�N�Bh8�'m�.�*�$w>�G�����m�O�~��}�-Ju��v��]�C���c�����m�Y�H8U-A��9��V4���V2�RƔ��m#<��5���H��7nݕU4��S]͂}mQ#%����{cd�w����{��5Ft�(�+�w�@y��x�g���ݳ���	U�k���n��3����)��\[`E\e\Bׯ݌��_?������n0<jǎA�ϰ@�����ӕ��筐�Z�@�G�����Dg�ȩll� �}�~��p%.]��i�5����|*�%Ø©���=�P�dX��ϡ�e�#�ᢣ�pKy3�NП<+�L_�
�=GC<1��;	-Ɛ,�?��?pE�=}"�������+���#���[�+d���bur��t���z��(����Ӵ�V�6��5˼��{ŵ~*��By����Yھ�V<�F��o��TN�E	���8T�+�*F5��=�}�K��H������˷��F,�4Y���i�oK���LCW <|OIQ
R,K��Tf��2_|E�� �h�ܮ�X��}�0��5�=�R���3��%YW��g���Fc?Q��C�#4����c�����'I���u�@~\?'p���<Y��=��\�z[��<�p�{�Yv�T�d<����P\̋ ���"�[%��E^�r�7|�����	 =��+��o���}�ʃ3h:iM9����Ry�:^uҼw���D���W��_�.�J���nDwG[���e��tuxq�.��l��Þ�cu�}J��|�1��.��KWcx�^ܸ9#wJ˧��^Rs44�$w�'���y�g�)�A�֖�)*�JtH8�葀�ζ6g�O5u&\����Aks��x�<'�g�vC�S��q���f��EŻ�~��o��`�1���Tp|��@�����p���U4� !@�0Q���Ѧ����7by0!���QA��G�;�3������,�g)�)T��l�<��P�ܩj��c몈��_4B�7���=R��khP��N���uv���$�>�T���ĉc���D'�_y����SY ����.�0���8�y`V߼}� %S�T<��7�S��}8��N�����^q�ݹ��<��.Ơ�w )ʨ��<h�sy$h��$�X���3�����Њ>S�T��~6���������S���뚼�&e���Y/K�3����^�A���MhCĦ�+U��Yg_!�Q]##�=�����n�G^, ��tl&��S/�3��NO�>�N]s���Fɻ�;##~<Dp4.o����O^�G��z��(Tn��(<Y��԰��3��/�΋��k�o^�:E�%� J�l	%x�oJ��b�'^#���"���_����
��3Ŀ�<��|3¯��U��Td����� �֠L�M�/�"�Z����������\�%$��NDo���TzD>z�qT�y�ҵ�c�6������M�U�ꗁB3џ�V��gd�H��5�ZL~��&�ˇ�:	���m���T�`�fM�U��Tҙ89'F9�$P�Ox���0�Z�a^UY��Q���7ؑjx�n�9{>�d�{֨*m��q�"A�L��4)u$7?�3�# �UL)2��&��6��%�7�0"��Z5����^ ?��f�I�|��<\��>���1A
�T:Y�8�=i����ܦ; ����fT�b?]��}��_{=^>����A������3b~^�?��-��3�Ä���,ğ �h�>�|������M�GjCX�R�	P�r� ��CJY����Z(o|�K�"�ƽ5цFM��Pi<D��b�����MC�L�0������S�į�y/NL+'��=̆�V��G�w��@e����X�E�w��3~�	��IX� �M�Ș�Eq���|�9qBk�ӄɗ-����Gz[�s�xtY�SB�y�x2�M��$��Q[@�T���[K��Y	��o+o���]r�+ �_y��x���ܤÞ��lb�S�=�����㿀_q�2r�v�`ͲH��T
���Uݣ��E����3�>O!�!�q���>��v���[ÚE���>�Z:�W�?5�����0e]�	�*����emeI�܌��*x�XX�)3�A��ϐf����Oĝ���p|R _Mm���-�|�$�n-f�=T�[�Q~�A��%���[�w�bq����'|����)ſ�8e-�0����,�
��|)jg�^H����ʳ�^�탦O�H	�+����Bf����W    IEND�B`�PK   <�WW/m�DE! ! /   images/ba63f8f6-a854-4b7a-ba91-7c7ad061d88e.png @㿉PNG

   IHDR   �  �   �n   sRGB ���   gAMA  ���a   	pHYs  t  t�fx  ��IDATx^T�חlY�؇}�]dDz{����wWۙ�.a�ҋ� @$$�ki�Ek���zУ��D	%P"@���tO�TU{S�寿�}FFF�����[5'���9�|�۟��tmm�^^�y���ƃ��o}��X]݋��E\\D��_���y���Gw�y��E���DwwW\\F�DWtG�wwtu�.���7��Z'qz���_z/��c���q��'ǭ��kD��".��3�+�Sw�.>��˺2e���|����M��xx>�<J���K�����$ʓ�^<-�K�,��X�k����4�8��a�L�.�����7����R������k�Y�e�1a�|��e�8���ey�>K˳ܙ6�5-�=�Zx�Ǽ������uA�泚�˴$�y��Yo��;��𕶕�>��N`*�d���xx��s�Z6y��Ϩ����tC������w)��~�*{9N �K�ɞ�����.���~�9i���N�4��\)���/���c�R���(�����8j�#�12�CC=����ãx�����O�����ڸl5w��Wǯ~����o���V�L�1H���10З@��F�0�8:>��@��G����ɵ���z����'�,	pzzhi%���?��W�o��/���.�OZѤ�֩��#D��dD�7"�[�p�xA�`�<�\v�u%!��w�0g"��ٱvZa�d>N��tl����Z��B\�]�4fL�4=e%#��iJ�9Daz�S��0J��j=	O^y�W��Q�M�v�<8�o	�]4��>!NO|
oOy������O<%2� {�~�Qr��f�ɄA�d�҆�gY��rS��|���.`2�p��H�x�y&L��f�������a�ٽ/�P��}�j���o�������9�tE�
Z탶{��`������a#��6`�s��D�2�����18<�C#�C�P���y�����&�{#����!����������|���?��_�/�Ul�F�:3��1>^���8t�B��d����ȶ��'�锎���l��<����r|��nގ�]��>�,�<Yͼj�3:G�����a)m�K:Jj�.�K5>���&蔊���о������SBϻ���?G:fg�ς/�{�*�����&u:��"<3�f:�+��a���Ӂ���1�(ە)�Bp��|
��K����	�o�E�y	[I4�t�� �
��}��W�!��/��*L��$~�HaZے�qX��]�6/�G��X�d�����_i }M\�������`��2I҃�2�i(O���?j����Jߌ�V����.��zЂ}=��jE}��0� 4?5U�+Wf�V�Do<0<��٨��cb|�6cըP��_?8$]w�����1�A���?��;������?���󘝟�����0������
6�= �=�����t�h�ӴQ����/a�lhY���q��g��3�q�˻0�r5[0b�@�qvvV:#s�Q�n�݃Y�o��>$X/Jl��g���A��o�+�3ӵ�'Cj'�����4ʴvR&,Y�id>��:7<��LAЮ��ju	"�!�z�P�I��e����>Mc��F�a��0dk�/B��K�no���9a����(uuL�˴@�;�T⤇t����l�o�^��lg��H��L�mo�M9V���;˧���7�K	�!�x��I���R>�P�}�~ۛL�5�!J�N<�[:��i�/���)�6��h���IM�����$���<�<[���	ңx2���>��ᆨ�;(cp���Z����׿�U|����?<��řX�6S���������7��:��&"�tx&�St�vl3[cG�p�@2������{�^isWT�o���aA<��N�AL��U�i*XBJu:@�>GDS���C������f���!�"��׾PZ�Oƙi���y%�� j�S�=�3=�K���>�mX��ƧZ/a-RV��>a�`b�JZ�!��Q��>	����E�Xf��Db��T�l/��h�RWj!�P ��7=u'l�ܝ���%sqXF�3���%OI��|
�%��|�;���)��k��n�ix�th��KV��l\�c����]8�k�g:!��<t��L����i5�P��Qw���z�aN�A���_��*t2�����3��o.���{�����q�F���p6��iL�Vcpp0�7�::׮NFϷ�}��Q�����?F�'b�DbD�$�����4��#X?<L[���Ś��R�` �aJLE�.�&���3q��\<|� V��D�yT��>,"S�t�	��C�I������F^$��~�
����]��α,�m�/�C�(���F]��	I�v�gB&8��VۧG�Ι�¢F��Y(+C��d�s`ב�M|�z5k���̲l2��!�M߁!}^g��K�v�e���r�7�&����Sv�aO�O���>P��"��{��Y�#�˶ ��:5�z2��C��/������Dz�ؖ|���dbO��pɌ
	�x������G�89:�~�vk�c166�6o��N���+q����|=�|�z�͌���r<y����� �9��ÍhP��b9�<��)"L@%:uH�c*m�ΐښd�����Lurz̳>�V3Rn>�(1i�p�p2Yo����:??�;����:�jD͡B"D&/�� �������	�&fg۩���I�8���Er�Lf�qN �3�=��#P)�x�T ���_�I	Z3渤���n/�����g�QÝ'��5��L��9��>i_�O0�����1WL���J�J�$��Q��BCi~�IF/�z��L'�FO�JM���K,@���8k�:��k��D�E��64��k��3�q� {�N��~�QO,���2�1m;�/N��}�s/]��3��������M0-坟�P.}�Ba4������6��6kZ�@��/�P�)R#j����K�b��eX0���B���<UҼ���x�[�wa�u���@b^�*��8�>�F�ӳ�U���:$C��[�x�x=��G��f��f�6AH�\|�������ěo܊�KU�X���>�)�5��! �S�T�DJ��Ն��F�`�>j �H�g#8;�����-M��8L���EX9;GJ}:W�B���+g���ց��L��ϳ�o�"_3.e�� ����Y��w�^bJ8�'���Yr������d_��?Q i��I'k&+EZ�����Ns|b���Vf�2�G��A�8�I�ݿr������R��jT�"�M��[B���)|xK{0��7� ���-m��}`9j'��>�l�A7�Ǿ�z��Ӷ�%"��nG�-��C��:>�ϭ��8H�&q2�ߏ+d|AӰ��WT*�����ܓ��:2t��3�!����:��]%q��12���;����z�X6O.b{�(��2¢*qJ�c
<j��1�޺6�?3ח�b�)|Ԉ&6m�-��ogØG���(N���H�'-�%��iF*{i��	��(�#�����L%�t��|�7)�}\^�a2�ҌDŤ�x:�}��st��¸��7F9;�fVP�d^M���rX�'���9}�Fu�L�!����TQ�+�=-�TM��ppQ�%�)��`���aRI,�p
u�݊Je�+�*������dhN��
��/��9��L�Zm�}(�����C�$sp�F�J�rM8�W�R֗uv�>�/�?�ɞ�H\��O���<S�B�җQF�Q�ZI�WkK�M���'FF0w1����x�(6������?�ѿ��_�2����	�d�B��vǺʾ�ͧhm�C��v#M�c5��8j¡u����n���rln�P�A60+0':� m�K�g0���~�GBqy֍�P$��@�+���"�L$�������\B��f6��oǐ�����j[��j�R��e�o�5����S����	��\��e 	�s���6��Κ��:Ńy�~�ҖD�LC���i9K!��ߖS����N���Z�`-�|��Hʄ�6�1J��܋G�
Ӡmmk����Y�*@��m�ʂ_�n������lfK� 
n3��Y��&�f�O�cD��N��C�Sk�Y� nߗ�o���(3y�2��w�����'}=( ���az���i�����_����V����>�����Ɠ�G���?���}�����ů�	Z�Yp ����`�1�����$��l�Q�\DiR�O��`+>���q����p-�w6b��i�[�Ђ�qT��wE�>Gex$&'Ǣo��?������F+�7wcwkD[<QSPA��%5�S$َr_nӗ�Eky�~����t��
�������{�Ο��0ݑD#Lڵ2���֚�ҡ]�A����W�-�|�{df�=��?��"��n	-���t��yN�0�6>���n�M�f�b�s��E^��I��5��(�hj"M������-}&�x�|�"����uu
I�(�Sp;��Fۈ3q���Sf����V��J�����0��(�vP�����4�x>?77n����LTF�cg{+�W7R�/��_�������"6�w���/��]�p��u\*hQ<a�%��GKO�g�ݪGg\��Z:���ԍ-0�~z/�����������������w�����H�
�aJ�lY×���Q����{��8Z�qV���T���H5��?����$�P:m%'iq1(l�^'�D�����w���-����a��N�^������6�!T��	��v��	/o����J�/�i�S|^�f��S�7j7K���t�w�L".N��%���GX2-I��DK��*Mt�KH���_ց��C�^
�v�G�W؊�#O��� 8����`����/�z=?��zͫp*�f���ƫ���'\�R|�7�z����{`IMn��m~��5h���
*�}��0�M�����beyw�W�o��r3��S"L)+������� _�����ۉ-4��A��o^�31�M���昌>�@��4.��bk�;�?A�~�� ��^�N[ԊD��C%��q�|E�666H�*6��@OH���E2�=\�j})}���>=���D�� N��i���P[Ҷ��e�C���]:����N�v�L�}��\��UJk������h��5#dy���$�N=��)�$�S�������b��[�YW� <���=��S�9���	N���G��O�P
��֡L~=,����C��x$b��
L���Lϳ�˓�ą$}&!��l�m,m�/�S����ӿ�㔤������f!13S�ɩ����g�fuy+�60����W�R�ilbq֏�Ł����"�����b{k+v�w�ݶ�d-�g�'���H'类y�-
�;����	�i ,q�m�� ����SKJ����pdt8�a�*L4����11��A�~;=�1Zs�\)��$"�,�Q�/I-�_"��;�t'k���^���J��	�%�ޕz�]���g}V:�kIc+K��Lg�IpmX����B\���?���۷��`>𜥦�b}�|S��L�)��0��*���d�&�BH�������H����p��v��w28[�Ef���Re%L�>�D	(Ӗ6t0�#Ϭ��)�s51/J��Լ����,��"�,��-|�*������Y�wӲ��r�;(o�`�W�I�K�1>=�8�ݽF��[I� .}9#�G�''��9u(��9��;����;0�	.���A�!��H���؏��2��؝��^���P�:vs�+f�\�LSfdd4�ձ3�F�_ґY8�̎P�.0G���2��V�O��<Q��W.2�x,Z���M)g'S�&n� ЧIdO��e�(ηD,1X)�_:3g��+�%�$�������X��an�R�ͤ��0��d������,�M��!��ءZ!��okҜ�LP;0��x�"$�|���g2��n}>�?p�_ybA�	s�Q���S�mC�tE;�z;, H�2w��W�͓��¢�����{�vO_�w�JP{b�:�c�'۾|Ю²��|��{�:�XX���U��=؄qNcb�3՘�����X]���!i�PN������4	�p?�w�����T<�*LR�#�����(���<�˟<ڎ���h5�X9sw;�h3gU��ęcE6��L����52�KMT�Q ��N!WA i���*D�dp ��/�-Q�M��D#¸�iQ����;�#�ӣM@�� ��W���n)�k兂�P���\���J9
�::�(JZJ�Wa}�4*.��2�e�aH�f�,eGx��&���v>O	KH
�m�<}�]�c����Ŕd\MS���?�G�)wO���h�n��}��nO�l1��m R�"�Ժ(��)�g�|�G�}>̶�җ��<(���D�@c�JF3EVS* ���G�XW�o����t�΍B�����&s�N4�CY=15Y���
�[3r'v6����v�D�w걹�s>�'e�d�l��
grvK��S���ҺG�9ӑA�[]��҈��}��
�Uf;:D=��%�Uk8�q��!U��@�΢���ҹ�2[p<�~=t�g����<�{G��cʰ3�e��Ι�jҥ�LX{A�̑N�����9tN�<��A��ݲ��`��-�4%"(sHh���՗�s0ݠ�Q��U`���ss�拂�:�딴mn��5�T�;�#��8���)�
�_ ��o�M=ꚜ�"���x�)�y��T�������k�`K-�g�Q�M�h��_���P�"K�[� �,.O���}���4%=K�F�,^�+�r��������>!oF1����ym�7ҧ�g��y6$�����������Xm4�qYJ|�/�Vv�~x���(���?e����z�����v~6�g��Հ΅��v`��;=14:�B��!ܟZ��2��;��[g��B
���w$��b��^�n5�`{�P%i��gp=��- w�0�uԊ
�l|l<��X��=�{{����m8}�AO�z�	��X� �G��
��OC@�H҇����{Nq/�G��/�&be
ײ�=ˑ�۷����f��4[�+�>;1�<�<6�aw����������I@��<����.�-8��a��J/�Tڐ�,����2Ba��F_�@I�9vT�D)6Sd���rM��Z��>��=Z 
8�0U����s��S|u�$R8Q����v]��`"_r�pXw)2O�,��3�X�+¨��Y�>��FrE7iz(��+Z���(8��I�_���,<�����n��㻭��G���uz�f O�pz��D�[/.����M�Í�I��������wڅ�h���I+��u&�I�$5\wb7��@t7��pŵ1St�plo�p�9O`.�K�����Dmb2f��cn~��
1dđk:�mlI�>��N�q�Q"�t\MkGup�A���N)�c^l���)t"��J���;���7�����=���a5��4u�W�#^|�o�h��vIY@�<��ujI��)�z����%�ȭ����yx�8�I�]��ۺՌ2�)d��:��"�k)���[�Dg�Le����)}0I�>�4m�P��4	��8	X�s�'K��E�k߶qEQ�6b��;�٧�ɓ��}fZ6u c�n�E�s���������)����c�j>�eP���7R�ӫ�rS��5���8!#�ԌӋV�������\�f&�op8G�:1ӋWr���t��닱xe6ᡪ�rK�y�����$U*==������~��� �ߏ�ȳ�ё����]����}���cl��d���`�!>�w���z�G�A��*8�0��Xlm�ш�,�F�Y�8*��gG��-��I+�Q�)��#�L��C����^=R����@j���RY�/D_Δ��#�<�����W�E@����o׆�WISڢ}n:JxۄV~��@Y�eI��CH�n�M�r-y}�%πW��G�qBB̏B���B��d���o|.S�����x�۠�J�������	�K9$����d(̃�d��V����kP���S��m�y/O�p87t|ӮO8/`����Vj��88lq�29�a���}C����y�ãC0WwV�PJ���13?׮��i�qm�w�)8�ա���w߽�j��!&�E���L-�y)���h�1>Y���ӱ�T��+c1Z���jض�S����TH�q^�˹��m�aD�,W�����L�Ώ���*��œ��?(S�Ą�j#2��Ī��i�8�セ�P�q��d�V����-�
:*�nZ~s12i�a9��&����f��(��&�[���Ge<���S��t��0P�%,�����\�6U�X���  n	��ǣ����D�BX9����F�ȱ�<�����Ruӛ�����Lk�v'���čIK���e�	�:�J��m���;Ө	N]Ƅ@���ɴ6-�����6�r���c��a����F4a������c��!�#'�b�8W�X��@o}Q�w%����g�n�ц��
�U����l�?VW6�r�0`w�qt�3<�g�c|��f){LN��ظZ&hmEk=N�v��&��S�k��l�17W�驑�s����fe��3�5m�9��~���.�@� l!��D�L$�JP�O�� �N�f��6i���I"�#���|W�O�V��ypJK��z�+�2Y<CŔ,Һ��I5%��$b�Y�5��(S�t�yK���?K/m*�"E�l'�3	цة���BD�WP��簳�I�}�q�g��"�"#M��������?g���3�yi����Hq���0-�����v�?�=���4�-�Fy/jg�$sh!� ˰ݔ��f{VQr<5I�l/��D^�_R˸��j��3�Wy��4���?o���J\����5Y���>��2{��]ߍ�'���h9V�=�e���˱|w%V��8���&}P�L���޹�,y�	�Rt�a���>���V<y��z��mģ�뱵�H g�n �$�bkﺤE��io���{ɵ�<����ܭ�Q�h�};��6-�+H�c����_�Q�V�p���F�٩�'��]������N?Ij��r���;�ӫp�ڔ)��]��e��G&����LO���]
Y�LWB\`ɤ��$�}�P
^d��J�:���h��'c#M5M�B�T��mh���-'�Z0�f2���򾃧Lv�0�,�KR\O���y��5#���U�?ӓ����4����2 F6�b;s-�'o-3�����?:m�<�6V���*LE?no�s1>`��W��@Xo�Xoצ`��8:@x��`i�W��$} '�6*n�[Xb�;h�&f�q4����M�6|������yL��>r1�v	��dq�����p-��i8����s/��tuN��q�]%S��=H	)7���I�\Y�����_݋'�Wbwo?�q8�OV��ѱ�E�P�$�Di�i"B��}��M����3*�v����Ο`'��Lg��I@%�!���͍'G��?����[����Y
{��M�H�%^�����q��x�K�!8�[V�F�:�Sne6>��I�j(ڦ�W�'�\B~Z?8O�6��f"3ʌr���h�坿���1�-+�a���Y2G�Ĺ���}�'��KPLO�SړkM̻b��r����	7G��~'���-�&&�Q�0C=�w�9>f�^+�Ol.s$M#v0)��]�~�{aơ������C(��أL�궰+nrb,z^|��;�����:k.f���X8�dC�U�[�W[A�Fd��u|�������a�����x�eZi7��w#������wcse�Ɲc�r\�s��j��)�:H+f�L�`�9e��N�,]P��wF��t:�r��(E�%t�Ͱ|�i����yK��O�J�$�Nҧ)
����{UH$ID��r&��g)6Df�ῖ�9N�����M��]5�{w#f��G)#��?4E'�+n��ԥ��� ���3?ϒ`�w>f���16�
���"�Lh]%��ļL]�j�Ӝ%�m��j.��%����`��?��]n��/��>#��J���Z�gr;��8�vvL7��*s}����8��9��`?5�	���fhp8'U���pT����/#�����0X%�U�����w�ul���8q��5�@\�V�%+N㗹\��bK� �H蔘� F`F�8����I�*Q��D�`,\�������i0�qp �b~����;ho#
,%���F
u����#�Mm'x|3��3;�4E'&o���:�&k.�������JY���Ϥ7���~��lh2`���5�r)�ZR��]���ƲJ��ߔWrq��S�Ҿ,���M� ���*�����	��񑖆��RoB	��3�B�߾�FR�=yǝ�`���I��m��� (O�wޛ���i?�s��#}�*�^jH�3M_`(o��<�:��,�;�)Ow���f��˨6c�2X�e�`��e�`_�-oG}ץ\�(��D}�0�3E���)G^��]}��{��^�:���Q:=����z��2�q��Ш��d8_N���֦�E�}ܟg�?�$+��!����')]~.�����QLť\^`t�u܌����ݧ!�!���hޕ��ܷ;(_�LM�;� ����S:�\���� TQ���J���o�<�s��:�� r�G�w붧L`>�A�����цjy�ʪίɫ�h�	HyH�N��y�����;g=h������m8=2��yKe$�LK��3�D'�PHg�d�D̃lɐ��s�Ӂ�ץn.���:[X�o��Y4s�b��8��������5�>T0��XPd2;�ۂ�,�Qn8-�st��J½=P���Y.�JNQ���h��T+����sO�pLM���/��N��&ban��qrV�/�u��8=s ��q��ng��:G?�bq��H����G�tk�'Eow������4a�V�p�ވ�����֑o�|u:$W�h:?�5�%P���"�x'� p��-�5�Ω�q�v"��V��w���M��pA���_� �c�����0���~*\8��TJ��T�}��R�%��OXJ Hس��J0��UY�W5M�������O�\ɭ�gj �Ix��M>;���ei_�1MIW�f�>� w�%���=  '$��$bSv��}�sjG �¬�͉�jP~�\KR�}��@��v[<����]K,'L�8t�4� �ym�s�&i�V�����}�������-���=�zӧ?���\	/��pSR�rW�A�v|r*�]��o߈�}������^�ݿ�~���cb��}�Z�ӳp_��c��S��15?e;`�ĶΉ�B�~�0;
~ui1�����K/^���.���h��"6�ν��ۭ#Ic�]oG��peG%3�%��m��5�
��(!/?1y��D2n��+�F%��k�4sI����6�$�[�p�	���n�r�:C`�,Ӑ!%'E���#���,K@�q�i>�x����8���S�p#A�3��uYF�N-��5��;w�Y$r:��y�0�H���|����e�.��<şgjC��ǒ���V�=�XM#�rM�dPo��e��䚑Xτ�|�;Lfx扰&���΂6�_�y(��ȑL_
�6�U�A��߳.���{Ì�0ؑ���z3�V���kκ�`�_������L\�>���[�޷^�go�ĵ+ñ����m���/2���w��X\�Ʌ���s�>{�ނ[���K���|.}1Q���Eϱx��+1<�_~q?}.�e�;�i%������uyѝ��v�b�NMϣf�bce5C����=��ȥ�4�HB��� ���J3�I�i��V�f��,(��+�w>�r�	�O�7(Ф�@�>�eOl�ܣ�ur��[��-��M*#ʔg�4��0��� *D��,>�f�@�d�G�I"�V��Ė- ��t�J���ǫ3
����}^f*t�Z.���g�m��/���vi��nO!�D��|S�@���S���h`��{:��UC]bo7,��?qa�l3iŋ��Ŭ�?�e�颩�'�A��Kt򛸓�)G��T_��:�˫gw3�'Y�|�����h��r.�L��&�0�_X�W^���P�i�m=����8��ƽ�Qo4��'�ʨZ!���h�3Lz^~�;��{��9a��i����b�j�#0!{��ݯ��OFKC���D�P�1Z�d�D����v�JywFL���t�/L���Z��뱷�*�T���(�s�)R��&sW��E��v�ъI�;>���A���v:;�(Q�$���2:i��ߟ�m_B37?X�Z�l��>����-�r?J�L1˽ĩo 4���c6�ЮI��w�QtB��NS�H��әj�B�h����X�Z���Mk�RN��>O�ti��@I��5Mj;�\�U�p%���P�OJ�D7�S��n�`"�pI���Q��N�8w�"�¢��.˗i�����(0���ք�?-�*t^��f�w�`�C�q�w�[z�����Tu���Y|��?�~�����~v7��_���z4`i�DGc�����̤�65�;w�u�9��4�nT���Q˥Տsc�SL���o rPB퉑�a D�_�ՍN�����@U��f.������C�}n��P������b�������̑i��,'�L�O�-����Y4a&k��Y�l_9˾�t<�;��|O��,�yy/Hjz�_�v
������S�o߷���%��%��)3w�,�$qxj�F���Q�W0HD�'���3Ӛ�]^1�D�� m�C��pRg2ߴ<\E�&�0���J�l��- �����)�UN�l�B�?�"���ޮ7�!���������/�e�C~��Sh��vr��!��v�O9 =
��"�N�pޭ;f߽�8��/~�~��~�_<8�{����}4������*�w;�J�T���@��\^�������`;~��_Ə����'?�0~����Ͼ���:�]溰3���2���Z�U�98�����.���Hu4F�*N]�(�m�=vfJ%����"���������?�i��=�m�2�*��i"����%��y�(7)�<=L����g���I&�����Y����^�]��-�smi��Ц�<:D��q>����i��$���i�Ϥ���߼%qJ[��|�y
��>/Wݺ�P%_2a�d�ia.#t����*ZR�Q��*�U�o-�z���lOgU�y����:��nGX�W,g, +�n])�}dM���p�+��&.L��9j���a���97�?B3�����G��c�V�H��H��Xn��u�o-\�9�� ���契��L ӱ��)��C��#��{��O�o��?�������n���8����gэ���c�k::!rll8'L�+=�0:k?g%8#�coS_����&��E��y:�^�s�d�*��>e��I�o�:�"����(5y�ϯ��$&N�㦱>$H�F3���Ô���E���1��b�t$&g����q��/�/.\Ċ��e���)H��a�����P��ߦ�L��$�̓{��;�c��C��3ǚ�fj¢Ւ��^N�J\���;��/�^���퓩�Q���I)�˩EVY�x��� M]p�▪,'�Ǵ٘��R�8(~P;A����]�u!F�+xwf�/tjp���:\A2��E(8�@:�,�uԀØ�]F*a�.�8cdT+J��L��<<�����i�"���B����@K��D�Vkq��.Q�j��d,g2k{��� �ʠP�s/cj^�6�C8���a�L�x��3���q�Yi�C��=wI����|���g����|kg��MagJ�ؑ�s)�ҕ�0�V[H'�?�;�\�18qf�]���m��p�G�\ܨW�Qg�u�$󀏲��L#L�]2��Hv��
\�ҷ�m�ª�GjuU~�<Aʼ���s� ��%�|�_$Ӵa)���\aT�IS��PޕaT{���țpf��w��1ϲNa����׬�����ิ�w),tK����JP� Vˬ���IS|Xґ����Nrw6��
V����l�ȱ��a���0�گ/�a�MNN岙��4$Gb���4��j�Ө��fPBM������6L�s�֦���3X�p$*p�kt�� �U W29WL�p,ͨ�HN�x��)�9hd@�*h�H%���O��D�.5�ү����'�YN�	����*y��T��h2���fs�:Y��RS�gyf/�e]�p�g�r�q��"���|N�Rt��t�{�3��DTr�������v}��&��w	v�����H���|��<�_p��6yG2�픅 �&|F˕6lG��3���:ě��Ʀ0���-��ϒS�e�R�e"�i3`j`��t2��Mg+a��-��хI��䆤mE16��fl�l�ړ5��=E{c{�Y �1�*�A�YJ�29ΉN�0R?;;�4��D���n������Q������'�����>
3���/����IF!���ˑT��M��a&C��Q���'��P�n�u^霧]%���H/�6�q"W&�O�(��+:�cF�R8�p�����$����|���`��;+��8�4}�vNӔt�hҤ��c6���`>.&�:���,���J}%������p%�X;�.uA8��Ey� a��� 4W%�s	� ?e.��7������y�஌��0�`Z�ŏ��C��������b�����2�������h��N�Ͷ�m�o8]���N�J<|���.�����l��,:͈��I]O&Xn�э���Fs,��ۈ�k����a���'�k�D{��sB�_t�e:��3Fх�B�$�d�wZp�v�>��{��m�o�����N7P��5 tA�zzc�2~ix���<�4A[�J���|8�&�h����ںbm���\����>�������l&;�ݱJ��?��]v�ϑ�{a�h;R.�s��(b�$aG�f����#	��B&�y�N�)�}�(LI�O���i"%���M`EC(�b�%�y-��#�:y
�:y��!Nh�D}o�1�?�k�Hԛ}V?J��{a���YB�.��������;�/�ZE�ml���L�|�m����|O��T���^��w�f� #�:>_�F��8\wj�>|i�1E'���|�7�����XY��-[��8j����N,/���~=�}�m�c{k/�:19� )�Ն[�� ՙpZ����}�p���Gp0ӱ�4�y\��Tv�(�P�����nJb���	�r��Eh>�:3�,��J�25I�#��x�KI�r�<��Ckyz$�a
埈6/׎DL�S�����up��i�y�Ϋ�SsPF�
uI5��3S)��+�A��3Az������Z����E���)W�\�	�w�B��2�y?��rZ��s�5Ӕ�T~�#�[F�1�Y<>G2f�/3K�2��l�GI��KyZ�|��:Ҍ���ȴ
1q�.�מ9A�%�nI�?�I��O)P�>?�U�f٥\۝��vr���d�F�4r��m4ܪ�/�C�~��qvq4毎�H�3Wcbf:�GF�	<�����mMWevn,�,Mb��S�p���"�^9z ᮍ�������a A��_D��;'ѨG����\-5���ޕ�i�p��Ϊ�ĀTmܴ��T���BLzQ���������D�o۩��yTf�|ڙ0.�I9�t�i�vL!��3;7M?����O;0k�g�^�8 OJm'l�廼F�%���_��zy��N��(p�3�0/˥�'��PF��T�F��
�{���샼�.O_Y�X+p����sAK��3gZ�`Rdq��BGђ�u2o�i]0�3�x3�Jj�����/uLs��>����mJ�1���_ه�/ߙ��,�{��\�6l_���O�$a�4���3z�8k��ЙIC�G+Fj���HL�M����X�q%n��L�z�VN�����+7���ɨT�@we��Е�P��q}h��J&''P���u��x�7��[��7=����L����=0&��):���,����q��>x���'K-&&�UE�R����|�.{�������$܈O�j)q
}���épu��e�X�X�?	�N,�Ց�I�\���)Eg��uKy���m[�Ͼ&]VN��b @�8J���%$���pP*�e��V�?��g\�;W֞8�Xl�wir��dY����-��AR��Jx
����U�ey2}�)�2���!J��s����+�ʺ͟A&�.���9��;uZ嘦����[�˼Y��&-h+�,K�ǲ��A,���������6�`G��\ڢ��.�p�jƙ�TF��~7����Xq��� ��3�pn���2��z�y������U�u�R:��c�M-,���=o��Ɲ�'~߶E��
������j��O�8���x��+���bqq*�ܶ��M��L|����ܓ4Kʬ{rs��EwT'�(s,6�Wcmm�v/����N��H�p���v�R�zfg�$�i:D):Sj�ؔjJF�=������p������kJt�KG����0��{��{��4x�lO�x��t�q�)�8���O��l� ���b�8Dc� g;�ʙ�%��Q�dd��4�^���{
K�z�|_����]�-�y#>K{�y�V}-��KmmyY/H�m7���M�ĕ���-Sx�?>�i��^<�1��h�����
˳2���~�kz���ⷨ/bo�����#�0�{���sm�Q�3�q��s�n!��E�	�G��vȜ��al�gk�/pva���֜��λo�q��I��o�!�5W@k��%����A��N��5ZR̔\j�T)�l\�$�L	�$\�&��<�>�?��y�t��qܿ��͙�� ����;X*�]	7&sȈ"/od����)aO'��=%f�Bٝ�>)���j�IItIG��y
��?3�D��y��M�d-��}�M�y��r3!��.;��Y
�%��פ���nv��������r-g�8�[�[괝�ٽs�h��/DXlI���ϻ6�lwo_��t��M2�����ɽC5
?�઎��22_f/?
��¨��(.yEmZKxl��K�,�[౜��u��������9'��1=;�D���_��.��f.6^]Y��0F�F��wx�Zd�N:��Z�K'�7�8ح�>������"����(=尗�(�sL(��2�_�� ��N�j@���p0�7�ƌ��$�����Z\�6c��	2�aL��� �0���јE�;s���=���� �`Γ#;�g�V��A�p���%B[��9R��1uk���D��9�"��x'y�m�ő���,�:�ϟ���sQ�2�k��}�pm��[�&bɛEB)�-�]�o�/w��l�
>�B����ӿ�~�ɟ�ׯ/$.�+�J;I���1�������u�.J5���8G�혙>�zmP�42��
�sJ+��#�݀n��*2oZ��?���y�pZ�D�J���r2�Z�����6���_� ۝�O�/�:��u��
m���4�<�.e���`���C�_��~3z "���ƾ��X_YG3�Ge��猨V��>��Ӌ�h�.Hӌ�G����rFҭG����k����܏��e��QN�D(��p���~�^o��o.¡کnHq[���[153���%4�(���������poA �q��{���|��rA0�J$��I�L���-��2��@>�_�i����i^ǅ�(+͘�!�;fM2�Y��/���yd�֗�R��s�̓iJ�����w�{ۓ���yڮ7}�Ԙ��#����,�d�HT�:}����}7�gG���&��Lǭ����uLYF��.��h�d:����z
N�Q;��g�����w"�W��ay��A�
W��n]��_��&�Ǐ�Nɟ<e�9M�9
�J}>κ��6@x.�Oě���8���=��Y�aާ'� ~���iQ�G������¤Ψw����p?�`�
ʢ�;�'�s�"	�2^���<��0}�xK�'�;!�,TaZ:�J�z�B-���7�y���v�5��9<t~!�m�\%��<88B�Nvٶ�T����P_lä2��$�g���\;K�ШN}i��Yoܸu;�ߘ����xx�H":/��|jʴ�"�<��eB(�%���3���L�4�ͼ���١�t�*Q-��K�^�,�f��QP$��-���YuI�G���3;y}���	�gI�5�������0�d-R�}t�0���;��d5~�����W�
�!��аC��\Bp��8�&�k�&^;GF^�
�ePX_���R��Sq�U�H�� ���+��������_��^��[���~�@E��~N���6
�lc�h	s�����+��?��ߏ��g��{���-�=���$
�. ��N�i&f_a��sv����0� PZ���C�`�مW�������{zx�fp�O���C�}-�Rq{9?�9���\�GP��Tw8�b�\p�_�4�z�!����1�vp]��������zn���w�k��] �#�nJ25=S�0�H~𯫛j���8��D�)��R�&b����tN�Y��O�O�CX�����ͭ)�i��Y̍N��0S�å�a}�{�iB��<"�HL��r�!D%�ɐ��k��rɤ�_"��E]`9��1uz0�5�o9���ޏ`����>:�������f)Y*��{��:e��7�3�����ﳌ�O���[n���
�'��{W�������W�����W���;,M��_���4�-(�Q^!ؾ��xᅹx���1��495�u-n#�GЖ9$A^i�"��0��<mg�]���:G�ʞ�.(A�C|�שS�.cSq�	m���t~�%6U���ӵ�"�/���bq�Z,,,ŵ�%,�ɘ���.�~���%�*�s�������o?�V��!����O|�ɹ������c�i�����e<�����]�j �Q�g`m�������p���0W�!���̙!.�����/���l�1�@(�δ�A�$�@�%@��Ο�ү �(�츔th�4�(K���y��p����8+�Ԙ@�b)�u�Iݝ�b!�>:��e���Lw��ǉ���Kښڔ�OB�w���F�~�3�����M,b����*A���7�q��[q���� �?�L
q�~1�v�~�{0:�\�%��0����������@H|�	m���߹w�փxT �)���s�E�*�A��p�!r$9�N��.ʗ���|f����m�I�8��g��;�#2�!T��38z~Pq6Q��f��n�G�c��6Z�Aۦ�Зw�W�����f��H��GQ�k�ڨy������44P��񙘛��㋘�Uz�F�dFw������r�XZ��,����޸����u��lc_vu�
�`2���+�|�g�\�F6�9ĭ�{�:1~�)�a�������X���{�h� ��j,,M��+F����ϑ˘� S$�����'?��|'B��8}�鳯���$�$�����Q:�X2H�M��΁0�H#I�*� \�T�4�yaNӖS)DT���h�/�>s�sg���Җ�ϙ�t���{�_z�F�����~�v<���U[Ӥ�)����G3R��r��kc���]ޕ�h���N,H&UW��pz��=�iQ8>4?ӋP>���}����*�lb29ǟuv�g�:�R��Ͻw?��V\��
�"�N����>~�����_F�dVA���|	�
^�e
k֥��vp~a�	�'h1��@K���v�r|zS��$�H��G��j����24�N�`�zfgE��lf�������w6�wcu79>
X=h�Q^�����J��i:2����j�!7ơPi��k�Nr��iS�Q`���)Z�y�Y?���7��͙��h����/���a����H�b�3ˡ�YVb�%F�8W��q��Iv�eI��1"_��tx�:s��L�ya
��A�i��a$,uT���4MH���Ju)h�4l��nJ�J�ZLU���<��M%�	0��l#�������?ħ����!m������ʠ1>��$Nli�C��񷀑��SZ�L�o��Xr���#Yd>�7�X[�/����O��c|��^����Q=�kד��p�w��&"��و���������y<XoQxV�Ș�d���o����%}^am�oz�����%,nZz��.�FR�g��c�~��E����X�n�*����}������1ܟ��'�l�u�1Z�Lg���X�iZi=�������Ø�-˱��LE�qs&��۪����8�������1+��,��x�T�~p�/m:vօs<��)<�k�1=?�o����r<��U<�w?��G�D��C��D0�ӓ��\A� ]���xNg��j4�XR��M�b�D�5 �_���k:��U����s_ޙSb�g�v�S��z9�ԑ�S
�	�� M�u����òR�[��ǩ6�O�%�\����(z���$�t����xx�Aܻ�8v���bvY�e	�������[��$m��X�@NM�@��6�^�:�czW�'�7�vH��G���l�Ǘbu����+�B-]F�^g]�W	̥F�6R���y�}���ۋ�]>�Q9�O�3X��~�Ԅ�:�;�,�]�u�p�*�)���p�m�ctl(ut��������C��61�+�gf��{�y=�^��������E�~�������_�r�����G݃}�mC�ؘ�E��D�v��Ez��+�޷��	����f��mexߝ�@ ����k�]�:�<s%n�Z�9ƞ����3�u_}u/~����O���c;��E�̥2���[��Y��&��Խ8��Q�~�W�ʳÈj=���F�s�&��A�ޒj\��tʷ���S��V� $T�݅}���W�G��s�~�e����h�e�w�j!��S�8��N�D�huܓ�)7�����!N�Ǘ�7@[�hC����O��67�bey#��;����3R� �����p�\���"M?���Ӽg��NU2�	�	�������7��i�_܋�R�I�N �.?34�K�-/��/�֑'�y:Qܻ����>��W2�wr������0F7e���@�e��m�\�<2\A���}#�f�Q�g��7��|�V24����
(��R���á�Y�1����D��O�G׹k���=F�mb��wh�F�Gh?�/,~�{�O�|�[��q���:���5Aw����Q|�> ����l���H�
����-$w�J�Ĥ��sڿ�8{D@ݙx�[X������k�;4L��o�`�V�:�~�j���=@�Z��cձl��xu)��a$�Xdή�<�2 ��A�W�^!���"����;/f��c)�u���P����S�X�ctu|�p���s)�lF��4]�u��vc�[N�F�'rS��8��ОL
��Z�6A Ύ�� �d���Ｗ�����:u�e@�n.5��ک��	��sxE.��4���5�zH(Sj�.'�@�y�@t�O9��2�̈�t0�����_��у�/�p(�e(
�����v$n(��$;.5R)}=����&}��R�R��[�2�\�'�U"Θw�#��kL�	��SW���[6�H3g���?���W�A|��o�w[ۇ�s[!��y�3Ǖq��+��w_���Qf�c0%A�b�ɐ�gt0᮫��ɧ_Ɠ�=jD�����=��n�?7�j��D�C��lh�8���Of�scc5�H���n��q�ŜYO���f� R�N��jq2�WB4�Z"51�հ./q�b�ݥ/�x�Q�$�V�h0����	|��5Ҹ�H�N�h�YW�8�5�\!4�� �SR�iYw�9��BH$as?U�C[�l�G����Dj��r�45�ę����È�l�D��b@p*�j�X�S�$���HjnM�\fCZM�O0�;_�t���o�ȟc��M�\���9}l�[?)磺��d$\�R��I�����uw��6�o�N�"�$9�d�$�J�s��C:�z��dd�7>��
r됙ȩ�~�uA�c���B����فJ�Y]]�.Mt������bM�sws���<5lig+�p��]۞�EC�za2�)���ж�$Z[��Ұ�&�\&�Ϲ��C�R�2z���;w�(�.l<��Qǭ7����pw�W�G��q�H2�*A%�c:E�}��LLMG��p���Ҽ�m���S137N��0�Ќ-L;�6�Dկ�幦��+h�j���K$���tbqc�����ccc15=�Z̽H��~|~m�@����
X?�F@���E[��l�ċR�����~x�"�Dgx�HfMO�>����_榣p���)Ks��qH�r�Ѐ�.5:5�.�;6!��a�P���g	$�G�^�,Α��QҺ������<0Ysy>mu��Һ��������.[�K�j�AT=���ة}�K�l30�=�Ŭ�lDf�tq�[LKҥ�o�@�_"}EC0�̾��Pxk�k����+z���y(����/��/�f���@��Z�S|n��2Z�eU����@�L���EtqZ�f�Hm8w������0�A�&����>���U��r��8sz�)�n�'�ھ�����_}��n�s��n iH}��!L*��Ώ�m�`�Ai)+�Y�m�}�܋�"�'��)c ^x�jY:������������5��9�z��_b��p �s��:�1R��[＝k|�?zq%2삔�bU�KC 5����DЄ���n��%O���/ӫMıZIΕ�����JF��{~�T陑,m'��֥��w�МQ���{�nJGC����0��$	�<�_|�>��C�qE�C̎㔈R�im�Q%C�=���a������x�i.��A5Ĕ/�il�>�ڀ��3qj�[VJ�<�Z(�Ҕ���N�������KżT���2Y��Vf�H���0�}FZX6�U�Z��r�b>Q#yh�*\�'����pN�݃^fB��>2����*��pS��굲�R!Y?����z����к�S�x�`+vuaΛ����~�y0WL�eq�F�hj���s�6#�'���PY_��`���Xt����^~��ČJ��W�u�Dwa���=/�9U�j�V��dN�?���οy{6N[H�͓��q��X�*Fm��Q����x�g��8v�D��b�49�IXΞ��_x���O��	�}w��9�ǅ r��R��!��I��@��<�L@��e�bj��9�'U2��,�4.o(ӕ$2H�2�	��!wC��i4�,�$�,G¢^aˁS���rU8d�CSH	K�-G�V���o:�������X�e���o�֙y��i95i�7��Ҥ��h����;��.���x+^�oJ�P�d�d��-�Bi#��@�����ub����Gԕ��5�0��� ������D�ed�
,���W?F����"�K������98p`\ܖ�(�4S]O�X�������4-3z���B{M�LP�v�>�6�� �5}мn���n	f�9.�L�zw��b{g/�� WK��g���QJ����$'͔����>H���Q� $E3#��8j!�1w�P�����:��d���3���XF�X���x��7���n���\"pqڈ} ���C��Dz��d��?}Q?�o��zv{#6��W���*!"�,j���&�t��hY2�������#�-cZ%A!r:��#����Nkx_�2K��h3����OJy��ƨIb'�cZ4p��6����v֟�L[@�9˗����5���N�R���$`�Y�|W�Һ 6p������΀�>aJQ|��Q3I��'
�l�pq(T��
QC�m
p�����\���>�6��4E�60� �8|\J'?l��L8����Ό���c���,>ZM!����]��8Ax��1�z0��T��Π���At�sc9��������0y��C�����q���)@��:����ԕ3Lh��ή����_~�T~K1������9���2XRu_�5�;F-�l���>�@e(�a2�����s����ch�+=���t�v8~����}W�~f.g.�6��/� a=>�����n@{�����G�����|�j��MHKBbHK�{���,����h�(}��'_A��%H��3r$�ɐUj#:ԯ{H�N!���ځ�B��Ǚ�9RJs���a	=�G�vMXy/�)��p��:��^�X��6�ׄ����N�O��?�N��(aN��Z����)V`(��Q��X�Y��e�5��~�N��"_�E�����t9�P@�K$�eO&\�M���*�I?��w�˟ZSg����_�2�W$3�inm�D16:H����EX�OFmn1��'������,\_�n�dk/�G����ь�ЁC+������΄ʡ
����F��9���g?0���˷���w�q�E�<�44�tǋ�%�w��-Ȗ_-!��P�o`0gۏ���AB�V����姖�ފ�^{6�y�x����f�ǫ�^�+ӗ����x�i�n*�q��~���Q�y�O_���OMYZ�SE���ٹmiΞ��w+:�:=n����;o��:�e��-L٦+Xa���W�f.	����9�SK��ܜ%[_8��y'�;A�P�I^�����r���,?���י�.O�T��XD0�`����4cl�S��Y�LM�R&��{��S?���9��|o]��6?`��6�E�#�>��9B��ƞ�*���2"g���G�(�"�*��>�Th���K�5]���.�ȴ<N|]��"L��p���1mzp�a<~��[��G��S��n������i�����۷��g�o���z���1#<�{�r`N�C\�pԒs���t�o�a`*�#�v�u��f��/�pV�j��i6F0=;=���Ɲ��M4W�@��4���G���!
v`��;�Iٻ���Kt�o�$����u���;�ؽ�g�^����x�مx��L\�2�ȱ� �oe`���O�g_�D��'�;��z6�^��ё2F"<��a���:Q)�@�)�p��v	�k�)E5��/��v��w�֎�3[�-Q���S����,A�H��
dyԛ�4��v&1�ߪ=:�{	*��r��w�ُt�#sg�$M&�k�OB��p�
��V
��8�g]�S�H2�,1K\�ģ{wȸ^eJ�m���#��-B�:���R^i��B'�!E�¬0G	�Nj�{�L82I
�x�L�i���w���G� �{�Ų���&f�a��/��}��}c4����c�6Ǎ�X��0���B�l�m�g�|���]����si�7���Q�SQ�he(��b�OM��P%ӛ;Wit;⧶teh\��ť��y��߾����%/(�RŤ�c9�w<�o^����x�VU��kאa������;��/�#4�{�61Ͽ�3:�t��
�+A�����!T��?��A|��n�`�aB�`�������Ɣ�=��iD���"���-�n��ґ��Ǝ��4�|��g�I�����5�(aSr}�ǃ�)[&M�&��ǋ&��~
�IT�)~F1�J4QBno@G���@�,t��Z�M�壊0���5��Qw�����H��P�N��Pg����a.�K�
?��ZX�I�\e��H#CY�y
2�>Iۄ5�_�+<�/}�{�O9i�dʡ@T���Wh{D�A��7ec��\<u�_�e���޻0ٓ�O��`'���g?�����`�����^݊���<>Ex��dcQM-����Dx�6
v�5��ǽ9&fj'Z��aUU�RϽ�L�.����$�.��!}E�k4��gE&��bj��z2���� yڪ26��q��BFP��<:Q��J�����J�i4L�uэ;I'p�Q�W�������ş����h��ԕS�����1���P��F>��q�n�{�#��j#�-��t��	����Ǯ�ǋu;��gL��̤s7S�
q�$QA䒧������GY�9�ʖ!cY^ywȹ�e^���\c�1��h3M��-f��D�l�푭�n5�G�X;�`y*���2���40�|t(R����#`R� G!zA!茴�{�7ͭ�,IJ�lqi��BF��������:�����YLcc��;I���0prmZ�ہG�P멍5Ae&�Cm�Ńyet�.��@;��l��x��70ʤ�X��莹���+Ø�ǟn���y���č�T���<���"D1��ڵɘ��7&���o��2
@�8�.�쫍��������뷗�ƭ+�p���n�&F�#9�q;:�x����x��Ÿy{&�4h{}/��;5Q �8����8<8N�gx�2����ʁ�^��.� ?�D�{x�H�;i�%�=8��H#{�`މ��]�Ʌ��c�KĂdNM,�3��f�C�Rd#qP&�ti.�l%}�:�&�@VgӤ_����Q�[���9.s��:܍���� �2g+� C��S��!���S$�?�$sX&��R:8���Gn�F����ق�� $�}��n����)xd��4��D)3<���� p$A�%2unV������!,]���;8���]֓_���=��2��'�쮕�Z2�g�\�#t��(u�����4���I��'a�aR�d&M���*`)�2xg��`�9�4i�8�
�ۖ��A��~��LZ#��C��av�~��Z�+��X߆�1�7^폛7��{?x6���gcr|0��r�s����;�Źj�������^�[/M�y�>m�˵����}����#������B�����=Oo�J��tҢA j��n�WŅ0����D"�w��z1n8��x5��Obzz	1~6�3�T�����Ә�RK&�?���_�N|���;�W�͡]�bzՍO���@�D���d�n�r%M!5XN��$�����։V�C����*�%�YG��IpHR?f.��Z窹����$b��G]�+y�p볬��4�d�3�r�e��:i!>��,E���	�'�'�������.9O�rH"AJ���`��w�<�;þ����0��Ev,5iZ���Y�p8F�\��?��˦�H����«5����`�a��,��ѭ��րu��H�-D���_��ѣU�t�'���t?L~������P���~sm0�~�g=�XZ��g�a��bcc7�WWb�:��X�fl�!0��^ƣ�뙦wX=s-��6������������i���K?B�s�4���]B��������.Wi���W�������+�d�N�F3C�J9�Ƹ��̩CK��p��dG*�;�F\}��};�h�f����W����9$��1����NݎZ�����W������ң���~��D�Y���H"S�ᡴ.�����>�CK�N�-�i�dɘ���lz��+N����1ͣi�Ƕ%z���C`�� �������t�3�� fԍC-�ߒ�. �v��-|�D�7�S�&�+�ڐ��F��(7#��99Đ��o�O��F;`^��4�0����y����F~6x�&��L�QΊ�j�ˣ���2��Y�ğ~�s2{aT5�S�3Chq�8�/�u(dԞ�j�bzUE~7a'�0S�%5�(��������r��dۛq�������.��O653�p� O�q��"4�K�G����V���p������Ӷ�Xy�����A3�<܈G��ڊ{,�R�A��5P:���6����W���ꉩ�j�|��o�d{�Snָ��o5X���+t����r\`rj"}'g�;!Ӊ���cp�n��ZZW�:.i���0��X�5���u�a4W�=� n�^�G_}��$�<���z���J|��^<Yo������H^�l�ݛ�0:%�-H�^:O-��6Ad�e�>?�-U�F5f0Ý�%vM��9y�dH�vސ��4��Y�<���R{PO�Ӄ :i�GV3f "MD:�<��-&Z��h/��'�(\�S3+@�q	��Ej7�X�/�p�OA��HAd \'~�&k�e{v��r�V�2�LH;�~��h@��@��:g�{�r��::8)����rt�kW®�\�����z," �t���Di^�U'~�0-�l��z�ޣXY^������!��q5��xoܺ>� ���_w��ꓕx��q<��~�������d۬�c[u]ƧG3�n��9�+O��`*�a��9��Gz���ą�؅��1@����IY����������w��Z�BՈ&^���c���IB�)y07�ɮ�zvy3sc����0[�pk1��F��Tb��n�S�����'p�qܸ=c�A�wX*{ޝAć;0H�O���'Y���kq��[1�0�4i�A�|�9l�1�hrAP�nחN#~^����+i�P�h>��+��?d�fF����َ�1R�t�Q&D�d��P���wנ
�iBvz� ϸ�AjޥV&�;l�T5Y2"�D�ݣ�i��p�,[���ԒjY�ʥ?��d���X5<8�|�N9�\§}�� V��
�DUi ��t��c>�М��'n�
O2���d�d��f�Ey�,�Vk�?Ӛ����ĳ�'+,*�����m�K�@NW%���_��G�S,�/��,Z�q$�Q�n�dn�;^zf2���n����X��\��}C9o���[��Z�<��Һzk6�7b��:���6�ã�l����΢q��,��p-��s�d�y���
��1j��d��ud�P��9F�:�-"�H���L�s��c#9�Y�}o� Gı4�DGId�h��'���� ��8���s¯��O3d?SWn���H�9|�͜�lY.���J�"[��R:���j0�9�k2�/��Ҏ9?jb+{W��׭�����9�C����t��ZƎ�ydpC��h4�$�sǱ�0R��a"�H�"uZ���)�sm�-��A02�D��g�I��f٩�����s�q�\2N>-�A ���ԑ�=�3�@9�q�S�M(Gm��A`���� 3	Y�)�sN��oM���F��4�l�ӶZG�_Z��i[�.m��zl{BL��gP�>(�G$�AE��
�ݿ�8=t�t��?�΁\Uq�8��ˍx��(V6��5']�8�
�0� t���vͽӜmP�� ���&�[ �)4j�q�c�Ռ ��fh �Lz/+ۏ����Q\�����wV�w�gO�<�x��g��ul��9�j���p*Ɉ4���.js���86�@���al�����@���cW�B��C0��C���F� �����K�y�뱀�|��[���⣏>��ciq>�jUL���(��a��N�I��%;�v��i�H2g�CXs�y��-GF�D�l���'�*Ȏ�l��T{rZ�̒�b�Ln�E2R���s��S��)���c]VjH�=�e�(�wY����_9A����,ҽfяI-�  �&�e��C����Lb��t�8��4�� _2�Ӈ\�W������5�?m��ӱ8X6��]>b��L��Q^8��3l �9h�X�3R��0��;��a���Z� &{��Qlᓹ	���u/���r��t0Wj�q���b�ֳ����ų����%-�k4�; �(_ʼ�:Jb{{'Wh��oժ.��6r�{��+0@�06��F�nX�������w��G'q㙫�5F�&�`5�Z�����9w꿦�jYS���_}���FL�ρ��h�q�i�+�܊������܃h������ ����n��x��e�_� ����14�\^!�N����Y����X��AE<X��T��D���>��h|��u�mI	Mp`.�`j���I�R�C�~HR;K��)�\s�»[j ���d
;Cbsq�;��G$%�L�3�rX���4�2�!�Ah| ��\��'s���t�I�J-M��b�"��s�0�:��ԙW@8�J��4�Y4!Ln�6�o�e�K��a�/K����а{��! �b��$��f�zT:��IY��^ s�j�j�Ӟ�����j2��K��N;�?C�Αu<Ͼ?��a�2�������O~����'ƽ�_���nLj�����<��O~K7��v 66�b`��=�x���������8�1���\�KM89?Mhdcy3�0j(�!����y'��܈mܜ���\��P�/�L���`�>�<6c̹�����w\�
U7ٷ���D�RR���G��ۋ���Z\�Ya�NI���@e��FGҮ��$qU�c�V�����ߏw޹�ۙ]�V��W�cav<�V�c���FA\W|���xxo�|���H�m��?��ct��N�����Ի̈�p`� ���R󂞃�\q�$4�!2!T^��b�H'�9�Hp�zJU�-���!�)F��>�^	VB��73�KC�������e"+��8�*k��*o9N�֐�l���*�f>5��X!�S������RٌFW�B��H���3F8�㜵~�
��Z$�q~ ��̜B��L8��x�e�n����fğ�"�8�+��O�~p�u�@PRg�T�ӟ�����7�~w6A۪I��<�����
n�>�YG�W�֋�Ә���������r��2<:�����i��[�?y���q[�[!�,LDuj�g{����k����y��x��baa^��/�h9�W��O������:��5N�H.[7�K�%6��8]�6�`�|�{�g��hB��3�]�8�y�i)�h�()5�0��#�.��G��OF��/v�C�^�?����������6>���f�j)0�{�S��!��8P��fe��'�gS�s� ӽ���Q��8� ��I�#0��T"qe�KF並iFՎ�ϛudk�T#������\ޢ�'L���ĠD�t6HF��_9�؜�DS��5_�x9/WWS��K���1({ ��6Ğ3t,g�c��c�G��0
������귝j72pR&��E
����.�9��Qh8>�����Γt���C;K�Oa��y���N�C����1=�/!�Kp}ގ�Xݺ �e�ht�Waѡ���8Aw�͈h������۟�_����gk4ؾ�=4��^3��b��0+{��8��ތ�8Mg�l_:�2V돉1��;%'Y*��dX5n� O����v;�^	��l�5���[��Lǋ/=����vܾ>'p�1���;��銾��=�&�b`wk��fR!0ͫ�l�L���o�a�N�P����4���w�e$������#//��1�`*;R�#,��N������0]���߯#l��"�i�o�o���9���z��ݴ�s�Q���,�c{3Z	�v���rm�Bǃ� Xw�*�C�Mm�)Y��������l
g���&�CkAB����Dd{a6�B�,ZJ"4���$~#���HQ�o's���3��3��|��dp4�ٜ�f`�%%�Oq���}]�R�\�l_�&�[��P��2�t������~�$#�Ћ��H�k��~��t;��8���Oӄ	�S�����=E`XhN��]���ŧ����fl7�b���ѹ�>$��(�ј�����0~q���p��E�ZY�6���M\�u��"H�k�Y�7����`���2ԗ��;9#u�L'"��cth8g'�ͷ����ٸy�F�]sҕF�?Y��kg�W���3��JkC�uރ$��Ⱥ�a�p�v��D� ���r0Z����ՙq�y	�H�Di�a=u5a��&���{]�m�
2Y�$-$(�i+]r���~�Z��d!���~�ۻ��g�N�D�xr\NiEg��t�5th��`;X�T#�6�AI-�ep�ZZ.%Ҧw���� t?�����J�9Wն��AC�(ML��
ȓNS�=T�9�L�������|��l��!w���8x;�eb�CE�s�XQ�I}�5ڃ �n�S�!Hzȟf�Ie(�.��#�-`&��9	��Dr�: N��1JJ�Ч����:�L�e��-�=4��O�=���0U����i|.T��g�ꭅ���;�F�s\x�,��ﻌ��������_���������.�"d�_f_V^ >{JB���i[uQJ�-��;�qp�ᾘ���n���
�[v��Q�n@�1����x��I�on���nc��t�� DF�(�_#9��ԳK~����>�Ak���c�;����_6�j�_[R�����v���T�<N&�<oB@���NC�L�F�9K$�&*�!4i�q4׍q�i(xva:� �}��8�R�Y,�Dp[6�YQ�G)��k;^i����h�q>��'w���;G�����Ch�&�̣ʑ�J��BM��:�
@��a���#�Yܻ���fDȩO� @�nO�G�\ԧ�Qi�	�Z 56���1>q��0�L�=I�l����-�X�O�I�����ӑΰ���B'�	���R�ڗ9ք��!0�.�& ҆2��Ca��Z������7�.�cZ�?/�^ȵ�]ஊ��5Z�3�vh�m�ǧ�s�B�̏��ȴ�)0e���Ql�n��>�_��A����cem/�'R�~��b�;~����O�ַ޾������}g��B���E��3���Eۜ��O��X^mBH��#!G���bzv6Ü��ث}qui�NWR�ͅ����v����I#��[1^��ۦ��د������o�@��b��*�W����\��	�$�2%��o�j���gm���I�; �|��`�䑃��>��JMGڌVR�&���-�r:�t�gP�k�&A�h�G$��t-5��Q;�:�C���b����f �̘�)Wqhz�<[n��k�
#m�I`���U�����h��}�{���s	�b6@��x��i�Q�Z��M�6�MI��̫1Z&P�/���`�^ˡ��2�)E��X���Խ#�a��e��r�^4e���X�x��$TT�F�I�t�[4π\9����Obkkk��mmტX���|��X�����Mώ�3���l����V|��/P
k��usYš+��e�����U1AN��q�1�-�)LXZH�S��)��M�[o����N�r �vf��J������Ճ�����g�}�|����Lf�����:3�]�t��b�|:����W�Ԑ�H��Ra�s�|����g���4~��������7�$c��F��GƗ�=!�ոzm�1�54��^OB�TZ�����r|�v��<gl��@����	ahk+��T�7:�^�xxp����4�(!_��7T�Ԥ~�7Jj	�3���d5�K�S�qd$��d�2%	S��2�ug�F����V0X�p���0_2��K"KMf,d�A��L,��ft���ă&��I� �S(��ƴ��A�`~��ܙ�����@���jw�P���_O�pQN���G�����got	|�Mm�Z1�_~��-�W�������AFZ���v�i�����_������O}���q��� ���>1��N��~�ֹ��2���)__�6u�f�V��pV�L�[�`������]���bba"�ݜ�s5�D0� ����DU� � ���4��u�n\�I�:�n*�����k�w�17W�iL1�-Ǟ���i�0��A��12��o�Wk;�=22��	��[19��5C�0�8�"�K��ӹ�����{�ވn�&��3���r���Er��~�CO�he�?����/8z��� gs���ud��v�(�j�A:�H}�IFS%�P��&�i	��7<�A�9҅��8ߩ5��Θ���e'���U��H���}���_�{`��Ս���O��o�dN§\�\���xr~^2��A�4�8ru4�b_�KI�I*. �&�J���ZK���4�ik�J!`;����B�~��S�R�������'���(�޽��M��,��:�Ú���
��1�݃��9���4�2�ס�>��ȀR�0��kOv���$��VU'k9�C��1��x�� ������\��)�n�:���ꫯ�Y]���nU7��:�fT��jW%]T$R���m��T�n���L"Î�ze��'�
N���V��g��w��)C��Ov>Dh��u
�1H�����4�A�kKs����P"�ID�ŁT�z�%H�A$nbء:Y����J �!jc)���xP�u�7��C�S:I�:�[���]���<R�F��Y���S0e��XmW���.�`t��ȫ�D��7]Β������D�_d�5<�X��eZ@x,c;������׺���0$.��n��"M?�%�)�K�5� �k�����eN5�X�X�aĲ0��*��ɉߌV:� �e����	���vq(��`.>B��1p��+u
oWW4��q�0��u�/�G���=c%H���>%C
�\'b��v���x�����D"ji���zǴt&�QC��M��3W�����@��!n�a�8�1��F����!zۗ���bGF���t��+g;�8WO;����e�Q����,�c
��
U��W���z��.&���88��W�}7^{��\K695��.,���/��N͑@������J����3�|�`�K4�	�O��|����%v��L!`��g�V�~P�4��.t�Qō��OJ���T��Γ���).�w�S�{:8����`4�>�,MiNm#��N4��#K�[�#Lr�c�n��R�z�N��r�.�xQ0�Ӹ>O��h]��ޞ�:b�rS��9`�����~�Kр�}��W>e�$�/�c�`����y�j4T�(n�g�Z>.�ܪ�1D�����[~@�ȴ�`�\@k�cMhZ��Bk�h�����0��Oqgp��6n��ى�x�����s/ċ��/��\N���%�֓���ŃS��{P6.���/���W:ьw�E�:�O��H�S����ͤ&gF��[�~����*Ʉ�ޅU�����X�{d�&sv�=f��;�S�PCp�����0ȃ0k�#G���i�ݿ����w_�w��z��Ϋ��[��3K�����x���X\�����싯�H�y<�{9���	l�| sh�~��	��%rvĸ��E�'�q��I�t,!q���I��#2µ2�	�p�yܽJ�����12�>�܊�cڨ��v��i���f���c'4�"��b�Ӂ����J��=L	�	��	j�g�akb��~$mc�h ��R|3��������a F��������a`�:�6�y?�;I|���&��5�Fh���HdS��>�7�� ��?�/�cyyx�I�u�9~�0��}}�i��d�Mn��:X�F�8'&����G��w�X4�&L�n{m[vw�ﰌ�׸��yZ ��N�r�܍�4�e^5ȣ������l+דi����LOt����~�����η_�k�g���^A��/<{5�����m�ܻ����ߦ��}�{1;3;����n��M��֥��RR@��'�_X���Bfjf��+3E[�$JONұ�9�dd�_�Zms�9l��Jy��n�zm,�+��� L"ǐ�h/�Fw��ķ�5�[��ⵗ�$�LqNƫ/���/,�l����h���G����0��/tL?��>{~��D�6h1}��@������jP��(]��4R�sPG3��Aт9N�6� F�05�f�#�2exkh�s���n'��TV��c�������jR+d�Ab�V+113�����=*`<�\���`�ζ� (	��Q"{Ch�Q��1¬N���w�9��-�X2�_�<&��_m��nھ>�I$�K�O�\��gV�ۺ�wh�~2�>L��1}�j5�{�L�@~�ܙ~Euaa6&�j�����=�|�!��j�7"�<���I��& }ҏգ�W�t�V��-���#�Z��P,]�Ü�B ��Лf|vxm2H���T���6;�@����e���b�Z����8�Y�������/j+>��u[9�f�k���w8��fc������S�ۀfX\g�6ǚ�
�;ua��ǵk3���!:��fU���	�KB�O7��-����39#Fmj"��rK,%�L��S��	��LVs< !¥�)N%ZȚ�;�<�49k�K�U�'+F
��#0��N�`@�������	���
)rt�ʧ����!x=�������d�}�� 3x���<Zٌ����[k%��Tj���Z��>� bee�p���13�T.H���!�N��h��V8#13[f'�8
Q-�!h��6�y���^��͍!=�/�N�P�O>9#��h�{ԹK�� S�F��j��Ao-�of�KW&r��¹��(�RLy���poLN8+c�Ĭ=�Dtf�!0Wx>��q�:��i�A�\���;i����۫�n/L@_�۟��ǘ�J�%��+S)��q%�A��'�Du̹����I��2L�����j����5)pi�&ǥ;��~���/�>}�Ϳ@p��˸{���R�Tp��p�|��7�c�����PC�xc:�?w%^~�U��<0?�2���U�'���+o?�|�E��C���1�0�v�[�)�Ո�А}}	*�r�֯��̎��l5�F�T0���w�s�B<���u$H7���z#J �_Fp�9�A���g�� �7��;?|+��A��+�)ہd�ӈh�����M�-��{E��@<W�wu=�������<ZD�-NS
B�j����v���E:���+gjw�co�O߃|���6#��+4s��p�%�X+ g���q3bs���4�<e2��^�M&�H�/��7��>t�n O%Z�������4;0�f��n���Կ�zѤ���Zp)��������
R��䧴����w�$Lly�'ܝ�ӯ9f���V���=A+���\KC���� F���t��f����d��h�u�eOW`����=�E�)��O���@��-&�2.L�h��<���H߹+MS���J^���>��~�� dסwg������]����pu*�����������1>3�P1��(����#�7{錯>����`^���5���1117nM����h7v�Vb�����^��w��Wk�����õ��s-�.�5�D�Q� �Ϗ�@�EL�M���48�H 5T}8��B%�����ʼ8%�Kp�n�POb�Ξp�jQ��9�N��M�J\j������>�@-�Ab�V~�/�2�i�uH2��m�$��ֵ��X~�kh���V�]+�sr����mq�A����C�n[~����\�2/�U�[�#~_\�n$)ֆ��mRh��\I^��.�L]��u����BǏʼ��_�:d���xMg��'H�j8�ߜ��J�̲Ϗ�p5�l���T(�������n�#Su�Q�:�e�v�3�i�@]�q|]#ʃ�SN�J��3�I��0鋩�7eb'ۖ��Q7�:�T\7��-�5�9�o699�BP��g��V�
Q��1O��j���66���t�
���.�	ں�������T��)��t���j��;���rC���H�=z�[5	��EI�{G���>��U��=ç}���}����4;�:���4�	<�B�4�ψM�`=����7P�]�v;[�`���[/����~o}��p{�Dn!{����seN��W3 ��K�,(ō�9&eG��|W���~��s���I���}�C��st%w]�I%�	M�=6I�O^'�g�ub=*'N�OT�j�L��2�az�z���'�J�8�gԭ����s�0�72���n���*��Dv�JsN������]���AW�	��ij+A"�A���������1
�u !���!��?4�m�38������a	#���������VZj='�a�N�U�|r��Y�^��Z�M�
�s2�C6�g�ǽ�j��/�
5�L�u}C��j�g��f;����)�:<�s35�����������b�H,�qQ���nѮXC����\YE�����J��?�2߽�7P.�нQS��6�5V���}���w���|��El�sL@?���d������ш���1���P�T���돌�g���+Ϡ�uƒqE�����юF�c������������S�U�	�����Sܫ���
Qp���5iR�j���_���GJ��8S�RLD9KsI�@�bR��`��w
_E)hİ�9vb�[M�_2����T�u#+13-C�u��e�JC�Es���d��F;'���I�b����i���AI$P'��l�����N^�N��(�y�x�ߢn�G�9Q�Z��F��|�r:�Zj#���!�;�T�h�8��0�e��l;��~-�fW ڌ&�=��s�W����7���t�ő{^:3�F�'�\���������[��_�q6a �X�P��_��'k�=��puP~��V�����Wf�D����Fz���RP���bskx/R�:��}Z-��a,���������Q�����n�[���_���f�XTn�ڢ?i�����o��@�(]ti�ȏ�p��w�4�ܐ�U�NQRJ��ԉ��|܀P�f�g�29�Ts��kqv0*��N;h/G�w�ss��������M��݋/�pc.�-�>�<67�pڗ��u���ܬ�������j0%���kƸ�O��J�Z;Y����k�����P���Ψ��9nC-��G305D�.3�]�?���ɬ�:�	D����duԙ	%^q+����O����8�B��w�<I�(���X�2ٸh�E�4~��OO"t���` }����,��W�ժ��D�2�`r��gZ���v���@�����v:@옩F���F��G�����鬠����"����$��Q��\� ű~��隠M�#���ql��?S䚱a���A5��k������
��ӀUm�P����bmm%QO��j��o6w��bq��x'N[{��h9���~��<>���⃟�:�׷��fU�8��6�cQE0)]<�XE��=�&� 4�v��a8;׀ga��"�3�ŏDhy��������sy��0䪉5�S�>�����O���À
ܮX�I�Z-^y�j,^��{c����������4�'?�(~��������^|y�0�]�ƞ���0̛.|>{`�7o^��7�G��=uP�bd8�#̂������O~;_�F"͈#Cü�m��,+�e��q��6"$��A�1g�´�+C��̏kLN� ��)G���9����NVc��B@pdӐ<��Mh@2|N�����~3j�U����Q� �&q�ُ�;�K��nS�j�[�!qU��Y�ULT��cr~�K	\>_���9��@�Y2���
W��[!�1}�:D�:F5�@p�@&���J��6�)�eD�L�S�wh�O�]�3N��8Vk�]�p��1����A�6�c�SWE3>y��OV��v���u��cw��E|}}��/�>�">�������x���?E�vtr3n
�| ����q�f���)c���4p�����sdx���E��s�8uV����؞��~��.���T��� �4~�R'�8ڗ�F5;�HBKiG�.o�i_���p��`R�B�}H�fJ��^�d?�S$�R�r��������A�k�
���W���������$L+�:�PGI�)�e�`�0�K	m�'��l��v%�	� ;iح�y�6r2�����!
5�KdF�|�dqx��s��2RFq�����(m�'Ѥ��J����3��ϝC0�$>���G�%N9ƩHN���ʨ,�m{t�����%l�놱e� ��ŋ�b���t����;wc�e��s,� ����Ԅ��3(m�K�t�2hDs��ec����v��ЂS�"���b�>4�R@�lBA���FaՊ�2ׯ�_'�c�������NST�h]=y��B|ggڢ��/����DzkA{����&�w�	�i��ꇻ�_���ɩx�h�)Lh��M��>��9
�(䆓W҄�<�ڣң�t!�X=���Ɲ��[q�0G&ư��bU]:� �+��Q�*�
J;�u6{�DN��K?H��/0>^CM+��bd|.F9��Keb:F�119��<���b���b\�2������b��9��]\�ɱW�^��@4X3FI##�͔��LJR����x
��f�B���n�pCqIH�Us����{���δ��S'4Q��u�U5��@)f]H�4����4��o�hL����D츢�2Ȱ���h�k�R�-
LH9������V�%+<#���	�0��k>9��h�m��(�(�\e���o�Ҍ�?5����������iPo���2L{|� v;w�VB����)�`Z��A�T�c�SZ`8�*dMOM�B��De�*�w��(@���X�Z��J���"��{�x5���-����E3��bfƭGbz~1^{��x��W��_��7�2���)���5��W6�p�����>�����cn~>�}��m$���W�P�I�ܽL���7=��d��t������<�U��]]�
���r��,�����>�;���$N�f���x� ��.�[��v|���㍷^��_}.��z<�<�Hx�F-^~y�į~q7��8@�F���Ļ��F�8?g�C v�D#�C/���|�dv2`��V��C���Vat�m;]�iG�VbЯ�������� X�ݒy{�uڨY���K������Fr?>�6�f����������5��ɚ���vq�p�m��ѹ�;�F�,L���Ś�d�=Q��BX���'>�*����l��NOb���r��ym�f����?9�.w��2��)�tA�`:��3l.\Vd}F-@����4�<����*�ԺF��n_h�Ԡ���}e�F���h�LZ�eപ�xx�I<��v��Ɯ\|�`��8�����ǟ��+�ҋ�t��;o���/�t������:�|eQ�(��ig�O�j7'h�}�������;)��$s#�3H��C��
�:H/tˍr�_ŴQ_�X*�h&��j۹��N��j-��8��G���@��<�N$;v0n^���޸ＶＲ�z%��5����n���9�i�XI%�;�3�PP��l ��Q��P������C1�73�&3�@�~P.�H��Hi���M��rq�$;�%����f~4`s� ǵ�Vvb��6�-$�3Z���)��W�K������~��O��dZ�\!P���|�o��sS`)<�pM�%�B̤��H"%�ϩE
�c���D��Dj*���}8�l��
�+���6]��>����	\e<Ө�~�8���5�O��.�l�R�n�y���~T�yX'.x�Y�5I�d0�1G������j�9�O��ۥ���I��SZ6-�\�G�# 禆s*��+��=����7��
�zkC��F`��pG6Mj����� ��8&�%̣'���tLϨ���
@'�AG�_���evkZhZ9�V��
w���h�� I��>��s���-�1��(��xG)V7L�]�S�VL�dgoZ��/b�ʭh��MH�(~R?�h�0%�J��i�!v�2���0��G�<��31�u�IM#��`����Z��Tk8�P�����|g`1:m��Ax��u�ɘ���126����H�=8���:�]��C��ѐ�2B�5�H�A_A��}Ǯ������ݲܓ���/�u�Ħ��$˒�d���<�L���O���,K T��F}�!��C��� u9�wl�A_Wm�R�*���rS�e]jug����0pj�V�cr�>QK	�&f�f����ZB��=���M1�;E��u|/Wӟ.��Ƽ�d2�LsNz�^��	p|��Y��(0�z�O��Ň��������O�7aL~LI'�oo����:J�(����E�.?���m�#pi��g#��	�H�k���`9��sxFu��ܩKAaD;�쀊� q:�ld�����t����x奫�w#��~�@I�	��Ӂ70������L2j�h0(�4$0܅�� �݆�V�5�ĥ����P��i�(�DZg*�fl�+\5����0��K�s135��H&�_�č>���aC����j��Q���pT�F�0�V�wŷfsMY��g���m>��D�����)N%�1��3bF�s�9d��
e�<<R�`.�Ԧ}H����7�B�|}�������I~�"�Ȓ�(C�;���i!����g;D�@q��~������I-��$E����٠��ǹ�(���Dbok[iDf�Q$H�OeH�i%�����};
�C��Ќ��2c�� pg��bu�w�#�҂�'\ӥ/.�9Ź�9�:����ܠ�������Gbc�/N�1��E0�C�`��6��2���/t!.jg��]^E}w#v�1Q����q��^Y��;��⧤:��]$#I2�N��v�ҿ6>�o���t٢X-"!�`������0�S��X��r��J �-0 �f���Kbl
��P�(�eI	@�J�R	Mbu>`N�"�~�>�~����_��M	]O�L�3ը��^��q��>N�Q>����%m֯�rlJm��C�S�c����-ѩ���2 ĩϡ��L-�Qt��ia�L"U2JN��q"ln�	���jxa�t2��ۜ)n,���?��̤9c�I��|���\�6�ڏYW�N�@f0a��8��\揖Ʌ���}�p!:c�E��OԉŴ4tmD� �H_e{�5eu�v��+#A�V(LҢ�*>�9�=��,l�p�S�l���I��Y����XYٌ�mW�c����4g�(�sB������t9�A=��	�>������l��B�#�G��yJ�[���,�������_Ń��g�<�1���f��
�/��P;J;��l��Vi���7x�l���v��.w5��X`�f�5�PjG�?ZǙ,�(�r�^�BvdvF����3�˖)e {!wA�Id���S+b�9m�%:�P8�ks �V+i��M$��,��jk	V	�l�K$s��ݷ�-���x�a�Q4����]���L%$�sǛJg�?�OD���n=9NG��M5���wb37�Ha@�$tHӪM����"�Jr�ų~;3'�B��E�a1Jٌ��A4��@Jy9�/��~A*�V��G�
��k�
��O�4,��5�71�vv��q�ށ	�԰��K_�j ���w�Na��߀�лp�};�WV���/��~/������WObmu!Y�n4�*�ùO�� �x���S��D�w޻�SX#�)�G�(�v��&g�D���m���b���~�O�S���s����O�㷿OV��
tI���.�'V2��Py�k�[o�~��@N2\|2XuI�:�~��E|�SC�ӏ>��G9ˍ>%.��Sj��W�:6"!+�Z<���/ߎ��I�F�阃��1�D�?�h-|�0~�7��~��� '&&���k�te?BE"���4N�-R����!��	S���)�!0`RM	2wt�2���߻v
��Mm����xNP�uj�$d�'Ӹg�IY�J3	I?�����J��\�40�ڣHm�����W�QeL�z�C�%	_��}�� 1�-~�F����)4%� 5م_���*	�r��DM�D�{��*opX���F�7���WSp��fXwgޢ�Y�O{��:9�E�$|@H��BWm�tx،��z�j��8lR'����ɉ񤱱���sp}u3VW֣Ѫ�H�|
I�׉S���?7n����F�����>\����~�O�=������Ұ�܈�B*Wg(��Y(���W��RK�}�\&�O�jw@�[o�qgeu'zh�ƈ��tP�O�~��WH�=������؇i��45��nT35e���oT,fE�P�ح�8 	��A�������q��O����y����d��m:��Ӄdjj2������r��@d�i�%'�b*�S��Ҷ�l8�)9��D����ãRqk���ײܻs��9�~��@��� }!MH�$�C�hD�l���tL�0BJy�op¼��"�2ez�V"t:������D�K�1(�H�����,��IB������4+e*�0�Ya$��0�8��gc�ϼE�ڗ&H�������k��(ۭ�u���2�Pƶ?�QY��Г��5�֑�l5Ns����Z�onav&^��X5���3z�ׅ�9 wH���$�v ����6Z�lȔ�PL���A�� ��9�/�_������A�Տ>�����QB�
۳S�>�����4m�~��|5]i��S1�Ł��y]��1�8�����.?��A�\�9�pZM�퇳��[)Tw���ģp�h���%�!8�P����zc�t��� <�����\c�� �Q��)�������� ��*d�/��b�~�v���cl�mlй�l��\,K�S#97P���d@%g���t�a�2pK�cZ��k琒�}h^~wC������댗b�	�0�Th�~�D��T�e��׌s�[��6�Nw�J%l�yɜe]\���#��\�(��Y�ܠB��1`�!�&�S�\9�FU��V�<�P�h�cTjG pU2|n
���ɩ��`ҟLe	$5�R���)���yy{��2E����2�ieMm�Dƫ���I.�=v	����5�#"Θq�8���Q�'q��v��np���H1mI��O��������g������œ'��x��W=���qR��z�/�/�Aʧ����F.;��4��b5t��?S�3�t��� ;�2j��Dx�l.���ݏ�-LZ�D�֩��y�?g뼿�X�������c�FG���~*(*R�1P���T�KM��׫&�G �V�F��:u:/{�h�H���Г�8���B�`�iv<�`4�NSº��E�g��a���9�k�d��t��j��/��3�S��8�j3�?�ls}�� ��'�H��K­$/ڧ��Jf��+jo5`���e	A�f���2~� ��I/�d
�h,�S�����BJFI�[6L �d� '?�b�֫x�Ek	�Qf���^_��W�]�e�K�fd����UѥL�R[k�l��Ѳ�a/���6i�9맫R��'�a����M�S�i� ��}�Ѫ�E��w��z(� P(@Kj����� smm��&��A+l����8��9�w�h���Fub!h��H�43��~���r�;���^�EG��s��a��l�8���'����F٥��3X�o�qgkïƛ�<��D��5 �f�����=]���*N��)r%��v��#� ��Q���]��鹘�]��k�A�DF*�|u*���|���d�L�"���SD:r???Ә�W�A���(�����`�v�M��o�j�8�-��)aU���l�cx2��Iv�^Ue�iEKv"M^������\��S����O� �ħ)h�el��zX~Fwɗ�$tj&�"�YWgt��)���L�),2�F�u�:���Y��z
�p88�0�^�y���EZ�A��=#�����U��Z��%�|T���m�A1���1�s5ǣc.�Q�۪�Bs�Z5�̪ϣ�>;C�^*�n�ośx)�7��5���#�EΝ�]ޟRO1'��>��XU�13=W�݌_{=�{��x��gbqa1Z�����y�9�����B�d{�..����S�%�h�ħgWjN- W(�y՚�{h�������w6�v�`Nh=ő�ɂ�,��t�$ :G�yT���G}��Q�ƹtZRH����ao�������x��ֳ7���+q��B̏��s7+���Wbv�/~��WQ?FA`"~jr2�'��ɦc���V�g�rwLOs�fE�j��FM�c':��24�?A�v!��FɜL��#���{ &gj+�\@���_'�Y��,5���iN��;5[�`1�t�IY�{��m~%sn���o�QSLfU 8hm=���d&�e9	E�����}#��-	�ā����0���\ԃ�m�E��Qs��B�'%[]�w�G� ��N�B�J�#��( �,�3��J3Ek�P���G��V�����j�"���r!n�@����빛�;N��[N0LO;o]��ߏ�~�j���q�F���{�ƫ�ǋ�ߌ�Ks��h==\N�(q�֕��:uN�W��|�˶P7@�j�cJ��{�u|1Wa�����5Օ�_��dnCl�Yp$&�&��<��x��AS�D��T�1X�4@���ч�1u��v����f��Ʒ����s�t�H�͌�f���zl.?�6��<���1L�I0�6�� M�%���b��v��@b�4I �if�T�hO1!��mh|�}�����������1��-9��e�0�HғX[�BZ��\�c{�(vh��Ӭ(��v,��~�A:����Nv��<����#��-�t�&�����Nr��٭chG���(��[�-���Ě��eM����X���M���4����\&�`��$d�"et��~A���e��}g�\ ��L'�S�@��<�K:�a�
6M����7����(��ѿu<վ
��u��/}IW~M��:�>*��ը��%l�|�x&���6��@�y]��[�G��_����X{����RLNM%�(���O�˯���4����C��%�ފ�����\9a�܇��[���S@��{ïI)�i�~��DEs�-|�}�7�F���@��� 6j#�v���0�p�ڎQ:��?�n\�4'|�Kz�(�I�Q$���U�7_�a`F�H��i��P��M�:o5�����*��D���9?pa�b��ath	����Z��Ng;[��[R�ZA}�4���%�ފ��:���g�)�p�%\?��K�Ї)<4�?و��=L�~�CsA�n��BH�S�(�%j�B�u�&����ccU�$�k�_�>���ӻ�t&�A8N.D��� m�3�n[g0@�,�ɘ[��"�jey�����)��r?@�I�]U;+@r��ag�5�ya���eq[����l7���\2�a��g������Ch"p��x�����9�+`H���ZL�ˠ0���L�T-t#�)a(5W���*k%�~?�VjB�=\�Oס��dX5�s`e����������>~��_|VN�꭛��0�e���?y��kQL:E`�������!�]$���5�n�?&�,����\T��#-�&��	�}�p���]��r�Zlr~:^{���)�C�P�k��czlaۓ��Sn8::��`bz,���r:�Sd0{��q�
>���V�ZI�� F%�>_���k>]	_�JHJ=CۮR��M�v#��ږpN��p<�1f��h��<ڌ�=̂�E���znv"�W��w��D'�M��gx�F�K�.�����g��3��R�D'y }j��G�����&�(� :��܇�-���{���)5;U�j1n�f��n{�ګ&��4Ow��,�0�~	u�'li�:Z�)nSq�ffG���(;;�B��2��4m)�ɵ�oj���ť�>>ج�o��B��8G��t�)��A�X��Eh����p��0���R��������%�R�b)����mr���(�d
h"��h���20����Y�t��Z�w�j��&~��/b}��_�VzR���)i�Z_~������/�����AW��6W�^�mK1<0B�@S�nq�ʍs�<X��_=&?>V�Z.���n��#;�۝���Ak<��X�2��,�(W��s=����X�Q��輮>�|�/毌Ǎ�s�QC�An�Z0����_��ؿt��<�����q��WS38F�E��'Ҹ�=���tR���o)A�7���Fr*x����?>i�^���Dӗrcҁܷc"wQ��4�hO~������K�������錾NTlDB�>wNb	�:��}5�)$�V׈IP:�p�E.阨��_���
���RS�N�N'n� B�ǽ!�C�rZ�>L�Ԍ��s,ib��ּ�o@�.N�PLϳ��U�h�)���pTM[�epk �����:�dN�"G��m�]�Q����ډ��5��ͯ��i��iGS۵���@}�VU�:u���.m�9��j2��C IbV�W\��"�kT ��G�,�.��
+ۚ��^�h8�m�$tަ�5'�����J�za)��/D��wڝv�Mxf�/���Vm�e����׎t���;|��;P�����$D�{?;��*5���fFf|wqv�JW�y�������ˏ�D��V�����~�e��,nޜ�!e��4"I�2�,4D�\U���l�Z�.�	���hJz�6qf5)����IS$�[��e�A�f��7�����x��J2/c�� K!%�CJP�f�u�Ի8�FEsc�$j���	���k�J,�='��a,�p6���&��+,Frs�L�Î����&]"���t ���H�DY|IW�_�����H�����I�Z��d� "@ݿ��2�-�ȓ���΀N����ej�����j#�U�;޷���Ӫ\�0*{S�1i�U��Ψ5}��+�5ӧfM�23EM3��4�����Vp�H�Kh���P�z0��77=�t��H��!/�k�NDpP�yu��
W�+���hJg"P&���7u��\���Y����k�a��+���TSXg*��L��.L��XX����7e�*��bna2͹]������xx�	f���ձ,-�m��O����$��[H�-�����s������՗���R��$?љ�Xw2��A���j��xkf)2�A�;��>ǭ�hb��Ҏ��F�j�ΐ��}���`<4�Sl����!��H"�v���uG�;C����B\���Y9l��2�T	��0��5�1S����m4�f��!W1�(6�	�s3�h��d�
	\)�c}�����c�mƓ�;��j�i���:��R-"����p��E�^��t9�N�VO�$E�0�'5Gg��f������6�;��mв�)t��\�=R��P��$�m?��#Ǜ�'̗EO����:�� ���z��~��6R���z�v�'�����w����ǘ�k�у/1y�p����~g�(3J���2��H��0<�m�����~l�?���?[�_<F9=Hȝ���Y�@W�aU����;wv�<6P�\��g�;�%��fտ�	�S-���t9�6��7J0;�P)�\P�Ņ���1-�]�����|[������7�W�7��2>��oL!��q���6>>����!�nl���ɓ��HӴ|��OɅ"����p��2�xm	d;K'�CB���;��f�B�K$8�}:;}C_0��j�]Iߧ��铑����뗺��HVF��q>�F�\Yݎ�:LzY�h�`~����f�Dj�}� 8�`EL:�R�D�赵�x�x\�ӿu��S��	����ȚG
�m�-��bD��,�:tTcK�Ί�T��]� *�Ǡ�P藚ީe�N���p�q$\��ݖ�@�G'_[���#7"�\D������"ܧ ��=��+������Q�K��4�y��g��yww;>��a��/~��4����E�Ո~4,�DT\�g˨N�3jބ��V��?|��LN�B� \���L�Ey���������q�8���������t�2���Jn�̫p�Q)աW#V:}�8�H4������{����2>���?�C��g����;g3��p�Ob����qy���� �MO͢!a�):┹��4bJ-Eʪ����ZH'��8��@:�4?�[+;:�l� �(9ۂ?g�����1�۲QT2�ά��gg���3H�,���Nz��������=mgzg ` ��VbcwI�$�F����+�%% �`v���i請�We���g��;�rVz�����}���{�1�s���f�Px���C�k�!�}Wm�PY���ZVi�Tg���V�AS�����0�*
-�~�<Ptk��0�W��5#~Iaa�
�pX%(�"*����h�Bó��B~}�3<4B�Y�ں�c�1����|��	+�5�nGI 3���eO�y�¼b����X�I���s��K��1���~6L_���^'��D9V��8�}3�?v2�W����U,I��WYl���g�G?�?��Xܺ�誘_܎%�H��kn�M��sx�A����$�W,�-�q>�%��	
D%b��V򑼮Bt[�t��ռ��g_�X����@����[0�M~Un��X�p���-~-��*Cc�d:Zg��H�u���h/k���hn��Ξh�XoT�=�#����Y�=�e5D��74���p��Ӓ)dy�&¤���]�cRȠT<�p&��Ϫ�&�nl�u�̽@/�[�(�1!����-�� WC$`���cpf�gb1�ΓF��3t��oa��]�Z^�1s�<F�W���f�Ok�i��x����fmBk.����ٴ��<hq-�p����ԷP�}�R�|7���}rɅ~=m�.�W�@�4��MF5*f��]G��):B铇i��WL+�7�g�X�i`Fp]��96-�S���҃e#r\t\fUA��i���r>4`��ٙ�D}c��~AM�g�of����'cmc�����fF��\_�I�emm7�1׷E}S7���5g_��F��rgZ`Wg;2И�fsu3�@�=�@�z�>��s������g��,�E|rIJ)�5Ͽ��k���`������\h�pV%��Y
��2��L`�X�f�19L���J��w{��	 �cE����0��.���x���x�J_t�����j�U7�~�|��)���Ǭbd����j��ӟbI���kH8�δf+����.����S�-|�US;ʨjL� ��6�CXi��45W��(|S�Q�L���<���j^O�_Yq�~�t�V�9&�ڮcp5τ���L������Y����|Y�p��I#�����,F��n�4@'�b.��l�c=B�=�UҪJ�I�(4��k�ku	h6�t�Fy~6t�JgXڍ�JQ��s����O~��0�6�td�O�<��[K,36���,
��.��B)wSq�Gy_��e�Oǃ3X�ux��;."o�}0���o����=O<y5�z�:*Y���Ӗ�P���L˹��8�`~���� ���
�pi����UX�h�* ���:Zg�汫W_�?!�c H��M��=%\͘e�x�>��A����F�EE-W�m��߅��z�}�������^y:�y�r<��Ÿp�d��0}�qz�1j4z����u3�MM)�҅O6::���t�<oج��e���Z
C�i-�a��N�}�����������Zl{��/C+�%Bg�ڏ���D&�f@ f��jZ_�8Ʌy�ͦ&� �'���@<>��YZ@�c)���a
O;��0���Lh<;��}j��M���Xܺ=.;r��.��>����>*����L�@9#�.=�oQ��R*�o�ږ�:�^^|̒�&<�[�,�Q��
���^��ܣ&����c1	W�"�蝾f.�@K<R��9��X���[$�%��*���bɬu��u }B�tW���@C�u���cO?_���ʥsq��������M~�Ba�q"���X^\�gU,�"U]|�lt�$?hHjp��1lZ_�f=|�D����6VlB[���殫�&m#�ŪU�-���p��+�=�0"f�X[��"����*ڱ'~�W��{�r\8����ɓ=q��`�=5��V�G�Ne�|�xS��51�����$4_g. �P �+�D�O���4>߁�=�+�0Q���8jۚ}s�d��Ɍ�J8�/�~�Uo�{�W��zȶ�Dp�Ss����,q�e"��η��O�c6�L+s�8zX��ձ��1���.cU��E����Q�ַ�5w���Z���sT
��,.l ��C_gf�cz�|��33���eآ�u����Q$�IBk��&���B}�3D2k��,X
�*x5Xg��R��C-OӢ�OG���F|�}E 䓩���JY�I���}�P d�b]J�*���\P�~�g&W(���5��n�:�v�G~57��|���{�3���	���u��4��{�WwWW?~,�|�8�,��o�iRY3n�AK�m�N^�[ش���H�L-�/�����#390�ܻ�@�3")rr�x��4~F��;Vo�_�B��8��s��64����A��(�=.o���4����7��~���,pW�s��m2i��t�i��t�ᬠu|�%�x����-��\�]]ZIGٰG*�oU'JZ�����ϯ�7m&\uNFIe������wo�}1����-̦����JiKH�����f�1�nl1&���y�vw[�)-���OΑdWP�;��`I����}���16��ǗcEgU�!�b7�:Y2�����U�O*�<���u
�Y"�]hԆ�.d6ri&��-k��h��*	�n�"&(���X��x��|�Fܳ��SxdŲ��H����&j:��b!R�8��߲��C�k���f�	�Ea�K�I��}�5��A���l�c��?D���O+m��R*!ƒgwC�L���������蹋�� �IG�6�,��Ę����N�n��:�7R+��\��k����x�����矊�!&tO��ͦ���w�,�L�Lo�A�v�ǅ��x���`,������caR`��-3�u���5�9P��p�l3vݎ�Ĕ�\��J�<C�p�;X�<h����I�_���vcf~=f� n�4|������V#�ØoP�����rܾ=w�L����.�q5��J��ϣ����#���!,O��'Mܩ�����hT|5��X�����N�R_�D4�sZ_i��?����eQ�����YH�ES�vZ㡑��t�\F�̮��̟l��*�΅d|_�����m��t���>�L���R�'p��ʲ,���̲�c���eIPH��=����ښ��*�LR�s��)%�JMx�R(ߗw.�O�~۱怺[����7Uofq����nZ;TDR�S�Q�2�z�55c�Ykxz*����AA�Ý�_x z���U�Z��ieU�\�V+U��5W�>��*�<֕_n�cf����p����^<�OtC���'�R�1<4=�v5^K�Z�ZX�@˶ �={�dt� LtBI��
���ڵ8w�����'��!@#1	�c�*����O�i"�y]�B�c�R��!��eJ5aF� �UG�љ~���ĄhmtӼ��|)�e�44T֞�vaY�k&�JZ����Bh!��T	IK�*-��SrRS�ˌ��w1j*��� ���%���2��(�1����iCQT`@��`�\�e�l4T��_ǎE3~���,�_l� �o�K��w���胔hM�����u�M�
F8��Q�{�ܠ6w�P&Mr?�����R�k�̍KV���p��B�\��ր9��a�]%����<l��kФ.�S��՚/]l����/���a�=؊���:1�����lQ���k������BFc��	���[׭F_�Z#(�:$ׯ߈��y�~�&㳗�݃�X�3��U�^YF��˴Hu�A^>����Zl�,�����{����Vz�1#>!<��u�����[�����<�v~��`ΙH��n'@��l��q�M� �+��w���B+m0:�6�L!�hMS+#\N��)w/{���\���m�b0��e�8\�*����^zW�,>�ju!���p���Y�ȉp�Y>Zjỹ���̣t�{5Em�[�;���:�Gw����9���S`��z'B�$2�S)�r=��-у�����l���q��A6!�)L��Q!V8<ڌ��ydnS�2����g��Tqz�tu�V�^��Br�����%i�[_�d��S`J4:y��|����`�����j� �LYw��K�E���<���EH�l�c�U`M
j�cg��K_y2}t�׉j�PzY�#-�V1�f�������0���}�����}<���Gq��dxd����|*��D�ɚG{�5OGl�!�7��1W��r^Z�����$c|)���9��Ŝ�X[qأq*8�0� ��.���u�0P��S�d���7|mM��ՙ8ܜ����X���޾�|�;�20F����u��`���\25xjc��ȍ��S@�Hxh�����=�gvn��2"mG�t�-UP�G񣲗H��3\|w��l���^�ה��z ��8Z�A�
�|	eh���-����%�T-%�fK������{�7j%���Ĥ��LeRfq��!�J������yW�@j�.�Ծ�E��'����#˭����O��x�`�M�F͎���»Ve_����az�%)D;* �v��L VQ{_y1(�N�2߹��������U?4Ӹ`z���p��$�9�ZMKcVNF5��u��Ǚ��ܗ�Ӎbmm����Z��N�{�~sK"����"s��(�<�wC�S���kA5��&�Hol�>�V�9��'�xjM�O?��ă�d>����{�U�I�r�D7Z�jqq+��pG� Q���0����؉���k�	��*57���@�������^L�݉��Ƈ�|?����[w���1�=���x����P�C� ��u� ���h��Nf$H�b%K��Ü����s�Ȓ��p�\T�'Ͷ �BU`��L�ZS��UB�:�:�.^CT��zY��J��ɐXU��C(�T>W���I�ӟM�x���$�	/
��#�`�e����dfo??򳤃8���fOK��`S��V"})�W����!VH�F)Ѩ����\��S��\��C	��%.�r\Bv�L�f�Z�I�;Ld�%�C?R_׭EB;:��<�%���Z:.����K'���}s,�'�ba�$5{�vY��ln�?39�3Kq�[�������x����7ߍ[w��6���2�'�5��L��\Μ�,���3��%�R�������}7i����zmvj�#(Ý٨P��~�P���݊9��s	�������ci��h��)n�t�J_ma~�܎�1@Kq���;�ӷ>�OoM���FL�GV�)���&���#tƱ��bt�[ɗ8�@���)6tG�vr�$�ʜ�SBd'ڶ��7ZS���Z;w�:-�c�	M��ߧ4ʄ��W���R(}� 
���'��2Oj6~JjE���?T՚jE-�]��,AN�p',��|�<J_ޤ�����m����S�kT8oe�f�(�Ң����LZ��u�A3*�M*\�0]F�Ro�t୥��xb���g*c����6]2��-1Zk��'�n���5ȜL���a�ZFS
$�
�kB?��g���0+�:���{Y���幗��2��gn�T��[�q��x��ٸv}	�e/�8��b���3���<����t�@)w'��|�|Ws͘kL����̱�vLS�-P�!j�}���ܘ���q�to�L�P��<j)O��$&ʗ��An{<x�B�.��W�Ѹ�6+�[���E'�����d�0��р����� ͇dp{�@-.|0���ޅ�v,�#d��a�тj5a���hSٷT��*�RS��je�*��T%�3����" 2R��k
�0Tb��v����dB'@�*\��m[H�g�J2��K�֗�xYn�`��;THH�VO�QW*���WZ?�9��d$�Ip�XY3�棚G��E�Q:�!�;�NAwq]!L���KQ"w�0�ŅE�&�Z_��y�A�T����n鍵���:~�E�zXh$��~�$���m[q�����(�!{����)_���]�������Bcim����	��L.�(��k�����u[(�����=����ȹ�c�Tt*�$Jq>=�r}Žf�vڒ�}q�3.���D~�S�w*t*Ɏܰǟzⵉ�Y:��e��!P�cAӄf];���sw2�`Zߠ?���S�*���I���/��Vc� Z:��X��OTA�[q���/��/�¹x���7�L!u���A�����;>'��c�$�2�`�Р\�T!0x�$3k�s��1�5� ����ɲ�����HV��~�7i=F'������Y�SK%�(@}���F�3�@2�Ѷy?7ڤP+�jGEH�(���3���uF����`~�s7�J5�\i��+\)B�i<+}�1����J���H��8�A�z�5j��f��b��?t6��O��O鬲u�ι��{�l���-}$���eD��Ͻ�(x����5����ʗE�b���V?P:�]�/1�۷Ƴޢ~�X���4;8X����he���t�܅x�������&��H*/���D
Gtr�5[�vU����c-j~}���H�57�tr-йt�[;���r)fwi+�y��I:���wK\�γ�C�F�1����", ��y|�WhA�S���X�ߋg_x1�����3�{,�~��x��'�'�FO�N�i����(�7���a3��3H+��OK�f	�2cdJ3o�Y0%k+����# �a��I��RAmŀr��&���
�¹��w���\�U��#�V,	�;�<C�/A���/"��G�h;�N�/�FfҺ%�z�"���h'�T�����dT��+5�׈d6a��8�*�&�w�QA_l�~�}�� +H����Lr�XE	^[�Q|$у�|���:������]�π�*�&e]����K�L��F�����m*�i�<+\~�<j�ǭ��ǟMj[�k�����������7��x<��鬐v�����q��p&��L���[�@.*n�8�7�}��18�&�o���o-o���C��N*�_W,��7�Eߜ�d��θ>�O���hl�B,����v6�O%^��PSĉ��q��鄖��lT���.ۄ	۞��%����슳�{����8u�'�z�cj�0>�d�	���2 ~�5Oa�r��T'�fP�?$�S���V�k]��b����	�6�dXB|��>�����[X��wby~%��I=�P(b=����{��v���E�`�������sC�Zf�|?�����ޑ�b�zx�!�jq3G.��e��='<a��ӎ���������Y�@2v�ܣ��j
&)M]�3A�1�h�Ke	��u�͊��2P ���b��I�5c�yQ���Y-��g����{v�mM���Ihl)5��V�AA���v�d���>�_a�s:
�;`ܶ�%��nt�5Ν����XB�<*yE�r��)=]m(�:�T�r]�Բ1��%���N"l�,���!�ynj����9���7����Uv�ؗ���H�V�(L�mk{[\z�\<���8q~ :z*�?��<r,Μ�L���h�C���t���pW�1��}4��z|���X���<s*���,`4��{���򃪎����[�G:ʺ
Nf�KH ӥ%��2������I���I�g�jA&v[��56+$R��l޷�7��m����SL�݌e�Euw�@,W���
}֓Aez���xv�n�̦0Hb?�{R�k��e`���őe4Z�4%j��=������s"Ӵ9Dv�Q���݇vZ��+hm����s-��k���	�y�Hl�\E�;��^+���|�kg5	�+y|V[�m���>��jiYv�g.���k���s�;Z�]sya�e1����z"{[nr��̉�7SG�0;jh���Co?��֢$��i�EG���{�w^����G���(Q�27.��r�F��U���3s13>�3����x�s��>���T+ �M��Be�J�D��N\EBKW&u�t%&dqf��'����T����/�BXz�`m0�F,�/$�5͞�U_w##�����m�U,�VFό�/��0ϽC�*�mC̔x&�GT�)_UtAڟjs�ҟ��H2B*�~W��d�=4��0=���X�DC�InG`zӹyw?o��v��SB<d`p�]}��=�ݝ��ͮ�4�a9Ip��	�e���P˳
s�m8Fր֌7�C������jB"�\�<Y�kjN
��ZZ+��ZTU#ؠ-��]x���upU�����%��1Nº�e����(�����C��)�v6d�����{����� >r� 
���3댌F��,�u��;N��ё����Bv�H� "2q����{�S�U(N�ªe�.�K�PQd4Vek?�/�B�Ҧ�,!8{��^]|��TL�1���ۃ�(�H� �x�EF57�� 2߷�ߍy�����݉���>��'��;������5K�vE{�QRP�s�d������O���3����ɘ��ː���sK1~.�K����Wh��ss<73�k\�`*Kk9	nz��l����̮p{�/�{n���&z?N�����x���;�_���~}��J{�<>��L��M�>3��S��0gy�dp�Q��ל	������t�7�7͘���VG��R��f�E`�0Jx�@����R2�@éd��2��UQ�����'��g�c+J�Ga���`��b0��BZ�)%���|�>i�����2�CO��5i� W�]��%�n��p�U��z��\������̦e݀C��57�h�9DXä�pu��,Ґi�͆�grs�����"`](�V��RQ2h��%���<ڳ�<|����3-�]|�ɉ�����Q��Sx�|_<�����lL�F� n���(�΂r�����񘘘L�p��|e����~�ZN�����R�.�c�������w�#Z+�XZ����6Z�r'uЎ�'̅�O6o��ʣW^��Z�j�����M�z���@�f�c�Eh}2&��}8њ�Ø�?�0��k
�p^X%qkbea#��͡�N��po2�L��r«c)Μ2�X�&�ǯ?��ѓ8��c���ҁ���J��<;^����$�$�epاo"� A%�9��wme�*B73܈��bU���R�n�|�0�	�-�P0��*
����u�Y���Q"�R	��iV�f�OM�`hL�^��� �7�M�����"�=��%���0�s'�b�	�yN�.�9&���f�ޙk�8���ļ�?30�H�a�Ύ���_�����7ې\KX\*�=���W`d��"�Fhh[$�y��5;U�EAˍ��`�?�"�}�.gdR��8|ޝ[
���cD?	��P�[��9�PW��p��J��޻[7��[wcs�M��#�N7aQ��)b�o�ϟʠ���b�zp���`��|i}x-���Y��͠EY�._�����*�`��yv�v���q��3)���5!�Y\��[n��И�SKvkr��w$�-�oj�ĥ+�c��~�r����u1�vgcmi�|+��h&D_[Z�F'����@;��`9üP����=���:���YO���ph�-K���X����ݙ��ɜ�9��d�dbh����@$��3 �K���I�,�B�#1}H�������,��Q�* 2��i�2��,%-t}<�edS���B��z�U)��?���#��8F���C�cZO���(�^+�j�x��/,���]$��(@+M�LKKk�g�/��K��		���^<����3�<��V��4�1���
��X�A~�B��Ƣ"���n����76�oh��`O�V��'OD�@/е+���1�Vx&''����
�-�`��,��y��n[W%���+� &���\��@��l-+'
0�c-�9������5��dKh����ap���=1�p��T#.)�aN�k�g �:�o��ZY��:B~W#g�fM*�fsu)ܽwo܎��w������ދ7~�A���[��;ӱ��SYU�'\S2��ر����B<��0>�R*�eMG?C\o���r�
��m1.x����N�Q�\&v�6�)��W*����*��h�
�d��Q�wL�PºͦD�R��++A�<����"�E�|�Q��أH|��B���c�_��`��Y�d;�Y���� �mb�Pվ����+E�*���g�ǽ
�Jµ"�����aP��ɭQ���֚g �TtM��b�U
��F$[;��t�l%���y����z��mӿ�V��g��%0S�� ޾S���E��%=�!���wg�rS�����Ə>�7��0>�v7>��Zc�-=�d]KJ._���l)�ζXE�̚m�Bql*���� ߳�z�΀�����jZٌ.�L��?���[��2����ՙ��^6�Ld��\�����VQȄ+��o��\�`'����[3ܺ��@G��iN�0�L��`���;�08�nn��k���քan���/}�%4�9�s�$�մ��3��[kZK���#t�il*��C"�V�h@��d�֭��@hJ����D���^�`����<�xK4��`!�WF4�Y�0D��-�Vj�e ��k�^ۆ������F8����9�E�;�A���x��F^Ư�u�v�������t��9��u.�?F����`%�ևya��?Tꗘ��
���&֟[Nt��(Z��Ŕ;��x���OE���Џ���j��(� '���,݌��vb�<�_=���X�i~����~��x��O���1��cC^e�0�Nt{�}����kbZV����h���눦�����ݻv3�'�bn~���������ci��ʹr���M-�oY��]ڱ��¾����r�v���_z!�U��']hv+GZ��PJ�e�ۺ���b��X_�F<ء�òX�]������L��!`N71�F��,@�Q�j~aP�Db)��0%j�yc[�(S��N�R��%�n�\i��	���q�)���. �G�H��H;�*�^�v�u��������t�=`�L','�}퓖$-�L�@
T���2E�]��?쏰�5'ŷ�K����Z_ѷ$���F�x*�a���e��IAH�K���N����ᅂ�W��R훰�4c�%�ɴ'ơEO���.>��B'����ڵU.K?��/Z,���Gsk�<�53��54T����gŒ*��'�T����
)6��VX�d���������\��P�]�k�����AD�Ys+]�7�">�|Հ�����tl.��?.dA ��4�R��$Fgg�W����ν�m��Ǎd� �Y�q{���gmnj	sk��at�]��FLek'���<�
������(v��#`ZFEz�f�Ԋ���&�oj�nZ�V�C'B�_���Ϳw>^��hn��������X_j��gO��p'�4�˧�Π����$�->���D��d(ZA�0:-SWGcb���hmŲڛ�.&N��^���"!�A��p�@AƇ�p��j��PC���<�F��y>���:�7s �ߝ�Yd�x��]�]D���MMM�<>�������؃���O?Ch�2
����D�6Ͽ]���S��j&6�Z����&���'�(A�昔X��W�ga�WkɴR�:�Syظ2��;a�7I�dh�1�=�뒋�3�:&M<�@c�OkŽʖcP��eK
s�|��U,-sA��P	�?��-�ctѵ67NZϿ(F�J�{k1�S���ť��_��_�o�����?�?�H,�����?��q|��E})Q�»E~R�Y����< [���"'F�3����$�s�I�*S�5�?~嵅��L���˿iI�Չ���Q�P���N��1s{(�����'+�_A@gu�	��-xu���+��_�{_������W^��>�d<����i��)�ù��5���ӱ����x��|/_<�%�b��d\��o�D���`�k'���U�wp�L�2��;3:�v�a֠�������R�Pv#�Z5_ֺ�d����&y���jU�i�PO__X�I+�O�65���N<��m#�zPZX��n�hD�����lN.����=�=���W;پ�Jی�%9?M3�+,%|��t �(g_|��
v��
-��J��S�S��΁���y��/PK�k���J��Lf�����gZk�	rG�!}�P��"�[�r�$�%��Z�-m��a?eh�����{w&cK�9VSH55��q�R_������W�x�G�h4N�9�Kmд��6��M���n��C�M�����-+�]'}������o�jt��
����ݑ�1��2�����$Z�����ф�騠��F�Q����@�M��`c?va�&�P��i*8�f�A�,`kCXޫ�T��d��j����V��>�[����!��yc>>�h6�%� #L��{U����Q�0D\x�`y,�6`!Ǚ�Š�F2�ys�kE<�4�~#�cM��p�Ӻ�lm�.�q�Z��L�i�'��FP��gYrO�O�Ǥg��)�Xl~��@�R"t[�S�O�OO��c2�b뵄��`ьԭb]�0֖��[�N����
��J67V�=D���/��-e�=Wkk%�U�.���9aqڀ ֩GY���_����F�f&�0	�)0��u�f~n9-�%�3�6�W<��]Y�����z��-��Qp������w������R�oOƍ���ߥ�կU�� ����
�Q_�C����|F���[Q��٪�Xx0F�����������o���A�E ��1rܢK��vU
ZO�S	07�Ύƥ���S��UI����E_��֒������*hӐ��e�53���=�(�{a50�y���j�g�|�cX_�h@�ԩ�{�:�5!,�=?��8VM��e1�驚㓮���M1�L�pA����uJz�{2���2�Mv��h/���t�/
�����<O�GY����bU<���o����ů1"&�tQ��4#,9�&D��
L__7��:�e���-�iqKƺ��h5����>QOwk�0QV��d�+f��2o���d���3�6�ن��A�b>�,�
�gllf^`%0!���V��-c��Hc�P�k��Ž��!x46�51���q�>�x+j��󬁱�3�l�P�u)w-+L��ګit���N��x��k{EW=�m7�xy��W�� K[�[�N1A3�P��V�e$8/���4����?������'?�ƦP2+)�.�'2x��`����o��tKDH*�: b3J�#�{0u#�y�[a���6(�w(�f ����J�Y�˗ap����kf#�<6�{"����ř�ChQͷPD��N�T�n__]�j&���v�z�p�\|�/��hp�0��G��vj�h�z��s���Q�YRP��z��Bc#��J���۽by��`���|���@�0�_�6)��ga����ֳ�1!+�>`-~#B���n��K���
}T��Q��F��&V�R�(�w�6�mhH�h���x}� H��*�2q
�(�pq}�G5�M�k��;������1nL�o:��
I.�Of�0O���i����7�g@k��a�m��󰴴"s䩧2��(k�i���F[̅�0�]v=�5I+�-�)D_��]�=@��D����sx��\����x/#��k(�,-�|������
cL���t�ag�*�zg,�g�Ԣ0U�.	��S`�9���]��eL۠�܉@;.C��Tf����~���2C�TX�C�Q�&����P�0ij<��Y���=j�ᡞ<���ّ�ßȨ4�{���R�iv�ڽ�y�~<�=3��1Z������i� ��U!���uq�T/�͚➫4�B%��5��c�6��"����,u���X#��?"�=��m.�=�gh�V�j!�v�r��Fbw1��tU���Ԣu�1��cIM��.���O���?T^r�ݹ݃�3��U`�L:1�w�I���˚�<ù3��v���
��v��K!����륯0��㬩�ږsjIq�"��_\e���M�a����1��9WW��>J�If���W�s�6��j�Qu���qI����kmS��n�*�tK:�����\�T�����R�4�`n#���k�]�Mjɡ�-�"���q�l���7�X�kY�-Q߂Bɸv�����6���pT,XD���B�<H�yv��o�����_�u�շ�_�8Vs!��o�T��a��I�'axT-��
�jҨ��6F�6�tr��-f"��M��	�a|�`�c��������x�g�b����0�����`������_�MJ%�礕gɰ~��2}pn:��-A|%.�oZA�V�c粂�$� ��m�`�qW���|,�������(���%h���!\]^�驹��
�s-$-U�ʤ�գ�nK�z�)5C
&��/���H�9�XpO����>�[࢑59&5��p��^����#���	��+V^�ގ����=k�{�0���{�Nr��k���'�6����@�t�WPE��pUdh�bkOz�
���dm���ND�W�1k���p�ڿ���Y�J�_�h�k���iѷ<,aim�0�Z�b� 0%���< ��O�}ym�_�Kfw���a���8��JK*c	�V����9g����m�k�MK��qw��da;;��_h  ��IDATo�y+�����r-��y� I*7���R(��y�8�������:�!�\ �piq!�߹W �cSs��-c�m����-������g���g. @���+'���-�ؐ���Ā������yvTk�~,�c��|�?{�� '�B��o�|&1��i�J�O-�ȹv���r
�Lin�kf�S����B�lۙ@�
˄,jZ���0��B���L�:�e����x9�X&U�]��`|S��6+)W�A'!���*1��أ����V+���]��
��Lz��o����G��x��8���<[+����r3���Ln������	��O������Ȟ��5�<]U:o��t(���Q��V6��ۅ�B2�$���4�z8�I�Ώu[\��2��|���`j)dn�N��BW�,߹4���/ŞD;ܯ���J��H���G?������~:�����[�4;O_���^�1x���X��]��ݺ9ܞK�@+0������艁hh�2��QU1�*�"q�t6(����)ڨy��'�Z��ΞJfr����Rl��{w�b��D<x0�|�I�o1@&_�m��5'�(����3:�2��"���!��˳1~�vܽy+n}v-���4>x����wމ������w�bu��n���P�\���eTgoǨ�U�Rn�W����Re��+�-��i��U�k��J�:d�31|-}�Tڑ�e8������BI�����u?��E�x�,~��-L?3��[��՛_XúB��f��*�p�u���A3��ā�0p#���iW��B��̮d࠯�ǽ�.��[����Z&�\_��<�޳�M(��]̥9،z�Rh�ۃ�����=��Ã�UbkXo�JDE���r�!VR��*����3sE�(
�� �*Y��gxz���9cqy+�[�2�z悴J��]s�U�?��-��,0�+(�t�ں*�?>����	��������N��{o��~�����>��`�,p�ڤ�G
�
�
	��߹#q��`~�na���UZ��T�(�s{�H�0j�>q����d�a�N�`�ڠOd���ߚ��M(�B%5�
�5���2�����.خ�}1곏��ǍOo�'�n���}o���x��O�\L-���^��6�>�OӯpX鷥�ϟ���n>���0!
}P��;��aR#}&�jQdDA!����.�1�*$��o6���A(��|5�t�b�~�V�dE P0�V�w�L��&S�Za���VA���#�<q�-w���	 p9Z��j5��94ȳ�`V���/S�6I�`;��5���D.�їX_��OO�4� f`��\Qx�oZ�}�Q���#���Sy���u��b�����-'Sy�~���ʹ�a�Чo��Rc�ec�nU�MS�Tl�V��f������L�XF�S��`�� �9�޺R Ʌ-B8��72�5-�M�9�w�|��d�쭱x�q���bX�.X'x@�څG,mg��� -�'��-��
�Sxa{���D��ȕv��_���
*�p�[5��k	�ݾ=��=�02cR�Z��a_ #���%�2?[�����7���kΡѺ�w�rp���`�8!��=}#����u����ۮ����?
�̞{�
�ֺX��3����[�����A��D!�A	����*Zg~f1��2��SX��t����&Y��N.��;[n�؇�aJ���r��M��{�r9����},���>O�(��Ϡ��N��ַ��(��)d��64�C?���Ad���rZ2'1�T(��Qh�=�<5����C|��p	�����G��:��Bf�{��z#��q���I7��� ���($.�����:��{�Ϭ���h���T�i%+��,
�
G��R�.ٸ����aoO�$|dn���վJ�Z�����4�UYxE�>
@��'_����2~�bM,�!4(�̓x�	x���C�V@Z��8A,������cᨰAM�nދ�������l�7��A��Iw���No��8��G/�61>�FЖW�A:�h˙�c�5�ANn���%6-��G�+1|jMݘ�i!(Q&,��7�uGGW_b�*V�P�#j��ճ�Z��s�1�q���dj�����gOk�z� 5��!i�@]��]��j�T*�)��Xy�����m�O&s�j���hfþ�Q沌�k(*��̨�76��'��,�#b��֙���J�"�kѝg-��l�b}}7����@⬰�Q��Y�E�4�"�>7��z�����Ȁ���R���,� �M���'0KE�ޚPV��A	v�v��K��aUU�]�|�p� �BW��� ! @<���0�bU慹fYe�@�v��,�y�� �����uS���4�����ee:�kY4��x/W���z��]��J�Le���N������~ם;c���\t�N��&,g��6�Z�є��=�T|��_��^y!{�J<�̓�ALLN�����8w���%�:��o�Z����ͤ�&��`�o��>�?M=��"˗�ح.X�KW.�6���Żr�~���q2��F���J�e�JR���1|�/bav.6�{zr���bQS���_��o�o��/�+�<�=�t������N�.�ɡ�8~�3vڷ��m���>�Atwv d��z���7%H!��Ѫ���sCUk�^F�	}I����=��D#�;h:<ƈ������pN+b���J���+]4B��qo�Pzaa��e.���.lk�j���
J��t;�{�L�2�`��)�I5��e	�lJ����f~���x09���"<�#3��j�L&�%�%��I��<�W���t�I3�,��lc��%S�V��qDP��b����s��h� �"-���k�-���d�F�
�����!V�!<�'=���x�>���-ю�؂?���QKY��'���OOȩ�@19o޸���am������SC�~����������K_,�z��T\�r9F������S�)nL50�q�l��ޔ0�ǲ��e�������J��(5�V|�F~���CiZ�k�?�'#�W�^y��y�L-��[��mG�P%�� F�R&KGЄ�*``c?5��C �'Z������[ѽ������#�N�ٳ}t��0	�8�X��_7�����{���O~:;�M�y�-|�Ա��^��L��[7њ�����^�OKF&
� \�k�dD1E�dDH:'N�вi5Lxb#����_.p���\a.ʸ2��U譝�Ok�uy��Po��Ӛ����^jc��r�Q܂��g#}�,~��Ȥ
�}���KjQ�����rp;����`�Ō�F`l����Љ��
2>��h���kH�mo�pǲ_���=�(]*'��<xQ��>���U� ��\A����N��z��[�L�����(|`.N��g�c��D�A�b��`��΍�Pȭ�'?޽=����Qpa���s����?/�p"�Qo�q7&g�����>�k��nޏ�n�b�<[z����>�+Ъ��{ z�e1��T:*G�5�M= �'�wB�.�i�}��a��\���K+L���j��"x�q��@x"��=&��W�0���Qg�s���с��Ǟ����Y;��%��
�m]#1=� ������p1O-�uPx%��Y)���G%����S4�{h�=�k�\f�A��6�J�� 
���$�*��/�=�ݝr��V�P��5����,�ae�nD�1��2�!�̄�2���[`Ԓ���O��5hjh�n���ݤ�m����pL�X&�W	H��z��"@--�|킑[+VC6X�����C-�a���µ������������W#�B�2�<�&oomD8,��a��-B����9�LƓ^js-�r��D�U�.xցj{�Kp�!H��H�xo��ί���Y�-�Z�X�����o���v?���o�s7�^n�u-k?fg΅��>����jBw�xW�s� ;�g.����oh(Z;;�6��CP�X^O� ���叔��cp��r$�)��������Ek�`4��v�Q�r��D|�ލ���X��J"�H��u$s���E|'���N��p73���*B��ގVljk�p�).�[ Ǥ���e�?�ΰnq�}�'^Fx�^97��	[D�!-�q�r-�6�������|LM-�	!,o�[	��c���HN��k[�/ �L��_KG�Z�՘�t��ZK����<�-����F���Z��˩?�P�����	�2� �M_�d�B_���庈�W3~��� ;H��\jե�p�m�Wl�P�
��z	�|9�e��v��g��G�A���sT(�;>KQ�Z��EnK�2��Y��3( )x� *�G*6�,�)=����㲿���U�R��li�5G0�9v�Eͷ�U��YW��k������>�٫˛q��d�L{\���iof��W���lܹ5�����JM�A<{�X\�t*N��c��b�d_�ud���Ɂx��s�σ��E�8�R���=��ﾲ�;7=��Y�ă�cfj!S����}M �v�7b�xXG%L��Xގ}J/�fg��7ލ�9x�V��O�����?hۢ���۟�S��c��J��
��ߊ�
L& ��ݶ�y�8�(�z㚕��h���֢He{y�3B�sk������^�'J����+~���Wa��,<�e}yij��D���G���M���;s�"���H��Q��'-��\&��L�ʸ#|o��0��$�m-��=͠(�!4��uD�RŖ��Z�|F�e���ii�-�ƩD�}F�|��W�]�%����̀DF<�߲u*��!�}B�XS!)Dy㟂&�J?����r��*R3�J�,�I������ �����G����PEIw�j��'�_��B�y�B��,߹oҢOV?�B��{�nd��ޝ�q��p)�j��\�Bsf��Wqu��X\^�y,���"�j��n�=8v.u�V�)�`���C���N�H����������6��Vd�n�͐��Z����>��0�%�[®F�@]\���w.@L�Uin]/N���D3篶Nx� �{�<2Z.�kq��z��z&������$/��ъo��Ց�vV�RU�9u�1<>����˫;`p�_<d�>��Lj�P1��VW�e�}��+B٤�>B�,�/ե��	�\��"O�T �s�T��O)�2�����/��d2}�FSaB��>7�*\̝�B�4�;�i��M(�^�W9X�Jxme`ɷQZw��e�]�����0.�[~��a���s�E@���8O�.:�8�|�-�u��_�,d�O^���צ�����*]�3���]ȷ�u�^��Q���?�lg[kn��@���)Q>�e��M��7s���z���r���eg��c}�M��Tܽ� >��F�����D���[�P����f��=�Lln��s��Oĉ��X���zƙ���Ԙ[�r�亓�?|�Z���p��iaa�kV��t=wXI���`�wgcq�n\�9�8��)ZO��7WqFe>>6])����%znч3��՚��is]�_Kk����A�01#��.�{���mQ�mioM�
� f0tZ:�A�i��T�l��S|;�ǳ<U3-����x^
���\KR0�&�t�p:1;t�"ʄXX˖'t��Q�����Fm8�{^����\~p{�+Z]+D��@x�c��s��l��vThf��ݭ�d0��В'�:�[
#��k�M����5N�;u7t�|ʌ��@���xK�.(̇A�L<�Ʈ��!�
��cQ:E���ʟKSi;��Jh.PG��Exk���'G�7�����#�R�R�G�n�!t��������E�&�PR%��Z�I�nj�s�gfq3P:������o**�=�^�!S�T4Ny����x�)��� �)%��G�"��fѼ���JLO�fh8ÓH�EA��bv|*&����fw�:ꝭ�x�g��'�G���n��Z���?���>��͍�?���韵vt𼖸x�L|����G�B=�0Ք�ܿ� -��.t��ˡtpFeP��p�WQ[����V�L"5�(Z#�Bj���r������t���������n�֑FN���f��|ZH!"HA̾��]�KZ).�2�f-�Q�窣M�3Q ���K�k3)+��b�"�/�b��*m9�rL�*�WR�\Z�7�Ҫ4�$�M����k̒
�gb�L���s\�O�׺�Y�"B�bau?��Z�,�C_ii?-6
Ġ2�t
��]�����ih���Ǉ�n_G�3����+�����p���U?}g6>�����R�N�`P85( �}M�}�k�G��Zf|ff&���ΥK(�R[��т�$a}�,&��Z[��w��?:���{4������=[*�����n��jD�%R2&U�91��1vg�	)�4L�0LX�v��F��Ls#M�T�e��Z-�88i�
&Xo��ҥ���j\�t�	p=i��or/���D���T'NK+v��t�i�u�]�D��Ɉ��]��':�	; �Dc����8N���Vs/5��K�Q�ey3�ә7�#�Еd���1^�/B������_B��xa�G����"S�����|82�ABF��`��o���o?M�Fv2��˞���<p�>��4ׇ�҃p�6�_�o��0�0���kT��bn�of�7Ǭ%�}���d5e���rmQp�Z���S)��)sǸVW��Z��H���_A�1s���v�ɖV����������cvftJ�F��������.�a5�T���1�EA-���:$)��s�m��3���7���cA4�Q�iķ4�Y�?��.��k�;�����0L(���Q��M�A�FԷj�^n�w�B�۫!�D� Z��c�dPw��ނ���	���GB* K��y�@�J���ہ���l ��.L���L�g����C���W���*Z�_�̤�l��>�31S�p(�
��C,��v"��,���H��¡���5�IV�eadH(���]���}�߈�������k}���c`3T���9�m��R���<�M���w�o97�n�PQh����5����D�I&��{��xt����r3��`l6f��YȦ�Y�_H�>:�R8�Y�_�޽L�а*�Ե��YZ^�P΅T2�0'@4.��k��.�<���0/t�w죻�}������-����$4GQ�8x�4�f��)s�Z�f9��Z�ɴ����q�9O��x���	|���%�C��P��q[o��� �M������b>�铙M����p1Z�p�� ���o���".m�'?Y�Z�����	�v*�k�C͕�W�|2�x`��)��4h-A�bl-B��������u���<���є�u�>&���/��CX��ǉS�c`�荎��8����W��^:�>3��i'֒ �>:�=��q�����nE��Èj�����@N�Z���Ț3"첐��z����-jqw�ι��I2� -�����0���||&��9���vj�cz��q�ص�B*_%�����n�X�u0�kc*�m|�qՅN#U
�$s�+��|��jSil��KY�y�����*M�K��(,>^��X��e|',�}�N��d9�NR=���f�|r},-�V���n(�o%(�1AE�͝�]J���U\&X�R@�\��P<����
]������}������V�tP8
�	�.f��u��"g_��[7��+ͤQi�EaҳҰN���p{�t�)|�����8w�,(�l���޽1��bA�^�c6L;µ+X�D=�Yiǅqw�.ϑ߼V�^+����;�J �swK͕G/���u+�席���[R�\4�y(�7�Z��b� L��D����Nf��ʓam7c*u~����_�r|��3O_��6o�r�9�ջ�q|�>ΟaP���'sQ��'�Ҭ[s�GNFow[��TQI�g-[�&Zϒn������Z:�N���*��i�2rʵ���榛{ dsn���I��5��M( Kʭ��f,(�fm�ΤU����N���h/ԛA0��N�V�Ln�����Id�.�g�pa����aq���Tqw���#��p��Zv�1�Ź�����+{�2[��:��|F��x�Y&�s��Vܭ-�� �V��>�*s���<��� ��G0��#�/�����&��Zf���H���.�+�y�G;'���y��ߴ+3��Tj�wWG�c���ߗJV����Ytǒzn&v�M�,�Ys��<����b��8v(�����G.����ͬ�~|+>��Z򛾭0S����6/�W��܄�6뇶�����	\$�7��|���p�n��~��WI`]q2��.e���N��i=� Nh:��KB��*#\%����-�M0�����f�j���I� DMc����Zv4FOWS �:[;c��F|��8�<̬Sb\��� [��!��rR�9�9)�#�U�q�&!/	g&�z`��5M�tw�с��ls�	��#tQ���7G_Os����"!��Zk�� 'Lf�~��<����Z����"��;HЯx<�{�`��hGq���ލpy�43��9-ģ"�	_[_��{2wRXRN�1��j���?���N>��߬���%�h��P\�%څn���u��7��TLjd�4�}}
���7��A��ݴ�Bl�e2}I3L*�����h⭹�>#�������
�}Ȓ�-f����.,-���5Cpt��4�e�ο�gB=��%��xCC�12RM�'o߉����h��iQd!�j��ʃy����Bi�W��S�U�Q� �s�©x����ܳ����t���.w�xQ��\ӮymFK��#�fr�~ބ8Y���)�imn��P+d�����V���V�}�14T�RH1�X���сn�1 fk�`��2�ǄQ�o !2�@��Z�O�/R��\)alK�{�F8���Q�7_�g9	����vw�Kvu�/6Ҷ	�L�f�x�!�����n��>� j�����`d2�x�1:2��2!��5�($��:s�Ff��!��0�Yii�Rq:�F*����g��� �]���@斏m����p?�:��-���b��S�����2~���<��Q�Qbk��{w��4�2�F���J������ctS�y��D��I�7��&��,Ѷr }��Z�d/��[�..k���y^@
�Z���������u��m0��BI�C��%2��"�P���,�:�B*]�g�P�������O�bsG�債i�ű����r�[��F�dR�"7�*�*���.<�Mh�b�6�7�삶�L�`ZhO�
JCF�|YJ@3�Z�x����㛿������J�;�	�F��9���([IWq��n� 55X�z� �0OD��y�.�I��F�ށ>HĠ<�@��{�x}Ea�	��0�L��-+�P��Ͼ��{�$��w���a����~
]�s�g
�چA}��U>��߭��ЄU(s�\��_0sdpd�n�djlAt���0�k�X�t;������haa��w׉ܲb�p��������B���"�7nX��w�&3Wv�G��jcx�$Ҙ��7�Z9�++��c������������#uU���sa='L����²
�����I?ӵ6��s��yQx��[��
�s�B�s�E~���.q�XYZ���P�gh�E*I����n�l�]��c��;�)=w�����ڈw>��$wc���^-��3��&?A;-<?OAuL��wآ�?�ү1�̗�����c�� G�U�λ2�k?˟�
-s��D�o�>V��pM��G��5�Sf=��8YVߵ�S�)ڽ��%Z�q�_y��C{9���5��U��H-�����{�-a��%!1�PA4�M� ���j"'ìl�[-L��5%��T�Y��$BG�H#lq�%��e�e�Q���g.��!�p�K���C�Ԫ���+O��9.j:�Yr�f샖y}����=Zn�Ț��N��a57�%�D��p�F\�,,v[
�@ػ�&czF���:��ͥ�OT��:9�=ŏ�ᙒ̀�������Z��	�M��P	�*�����ڞD������̪���H�?��3�Q�d�d i眻��ߪO�:��%�,�� ��<���e���o�\6`��TJ^�w~�ﶭ��a�=yM��B����*���k�ڊP<�� �s�%j��-�㣥�Z�Z:��?�o��w��?���Q`L��I՟���� �Vg�!H֘�xe B"o(�B�� U��.�����A�dn5��o������a,�90�/�|5����w�>���n�u�� N{u�Nlй=�K�$�>��dH0�r=�2��៩EN��Ǘ�I2�%��ҿ�dE"�'m��EJ���#M�1�)���{	�-Q�}���}��̔N���aB�0&N��Yr��r��G�tpa2���D�cYUe=�Jk1��������u���L��=�M��k�����*��ʦ.qʸ�j��x��-�F��Խ;������<��e�B�u�BKh 45�^�sM����E�;�c��l��2(��³eR#|
�
�(���s�r��90�C�%ĔQ�V�P��Mb]-��E��M�p���PD.���wYw̵@��9�%G�D� S����]����`/�)4�Jz6c0�I��$B���L��T�ČS�?���'V@$o�s;~�捸����_D١��Ma�8�X3V�0˻𻋊j;5�V3��:��U���p���y�Z>x�F,1m]e�"/��+Ʉ���ή�d2E�� k�6s����-��a��¸��}'>�5c!<)�e�%sa|o_SkA�\䅰j.C����p-iŵ�NZ�id����L��Lo� �<���I���6��*�n�!���tʅ\j�[���f���6 4�ON���c͋4YV�cEY}<O�&���`���
���<+!�S��Xբ�tykJ?`�?k�X_t�,D�;_G_�yH���x����wt�(�7��F�:�q+ �v���'�zrY��Q-�ӿ�m����I�-��A?j�jk=f&<�u>�
9x���|�Efv���,�:?����g�)Q�*��?�;�s_ ��#�@�	��sQ�#C�Z��%�SScu�����s�ș�X����۷cj�AL�ߏ���zk'"+�).W�0��z����&�>~&F��2����\9Q�\J2�oKTD��/�~5�=��k2�w����ft�ݽo�����Ïcb|2>��.fF�q�S���^��q��@���Jƴ>�b|�ᵸ��M�����z���Ń�w��g�Ʒ��?ş��������U�S��
2�hǩ3��3lm�����ӹ��1zXQ�O`0@��L����cսq�K�n��R ��X�ڮ[)�������Wvb2]���;:۴|>`5&3.�a�eڷb�j涵uVb����U���_B �ޞ�B����j��5�!�I�扔��i����5ZYdl0���-��0���m�լ�(3����naɅ�ͬ�1���@tˣ-�.,���&�z,��\yt��e~t����h�l�~�K� �6Xz��b�nn�Nn�=��x�M3>s�F�ڸ��9Ph�kg\+ԅ�����5W��"��p)ܞ���v�D&�tA��Ux&�j��J�5.�ߺ=�����s+9-��Z�e)�`1;>����Gߏ��7�c�������������[2nwp�N�V��k�s� 3c�mq���B����ROX��<��ךz_T4ҧ����>|�û�oC	���X���Yh�E����
���L��S!K�5��]��	'z�{���{q�Z���z�����1����N���h¢Q�X\��O�׾�R\8;3.2@�'�`��C�{S�0��%�ǀͰp�
�8��U���)�N��?	�:�OSW-�����.���N�=�|<ɬ
�di9���Rs��I�߻7�yj2��fe
�j�.���:.������8�D����j`\a���Z�����/noa���O�����&P��q�o��Z]
�U��6G]���+�KC��$�u��BVP ��X�l��,!�D��.c�ݴx���J�wB!т*4_��	�P*_th�C�f��̩�±�L�5z�^f��san[�������7��On�8V�����]#�F���v=	�vϹ؇��qPZE���NO-$?֣�3�YJ���ϛ��ng���w���]P� �AP�Ë��+�:]�[�e�o��o�����&�]ht����w5^G\(�Zv6�����]��6�x	]�k	�m2���vtv�����Rkttt%l�^�iG�ۃ�,¢v����)�@h�<1h��SW���b\�0��ZF�̬�=�� Tj;K��	)2������x]�"i��*��4T���I�aB�V�|��
�y�V:���w_��d�V쯖Wp�X�2��V�2�D�le{Zl���ln��#`���+�Ό^�̋�ւ�A�5�s��GZ^fa!�dRY�ܶ�-�����2����P惿�k�A�C��#rڣ�|����-+��8�\��7�3�ힼ���4���;���
x�]�g*i���lO:�T�P���S��#��5H��w����c�P��F��T�p���Eg� ��S�UD�-ŝ���ʊ�����}&V$4�����A>i���m�,{�s�2`g��]�~Y��6k.?z�I0��rcӂ�k�x`'}'�V�p�?����[2g�5'����GQ*	���>~�l�:{����N�ƙs}������3#��Ձ؁A�g7��IQ;��w�ر8���[�L5~�����Z�_�1&�|3f*��0��UN�p��֔9#��f��+��&r�UB���M`�]��1�]��� �������v3�)C��`E|_�hXiGA��J��V��}����(W��ch?�� �)c�n�ש�eZ{K���&ݪd-��FV��_�y��
s������u�s�>�K�%�۹O�G���J�R �a��Т0F.Ӷ��L��I;��&��tSK� �kr����x]���X��ghI��u]�⦳�W�ڤ�J��Cr[� .=2CC홖7r�L����䓏������0�z;��&���P8@}�xS�FO%2�^\lG����^;v�Wn�����iTX�����⥋���.C#E{yV���j����1����E!�f^�u�$�lQ�)��mM%oж�ֵū�~!�������g���q���h��X�����ܹ��k7��uns�u�btx a�n`�v�-�	!�0j$T��τ8	2e΀��El&�ҘH}��b%�����.
�S� 0�̑\E;2d��S��w�S�8Lh�����n��?Դ�r��}9R�˺$
��$dbI��Z3��θ�D�����
�!���Ȝ��\I� �N�־�L�Ǩ�	�)`<����4��'�0q٢M�[�ݼ�e�g_uɣ ��dΕ3� ����P!������M'W�R���
����GE`��
@z*������0��(�ē6���������ͷ�AY�����B<�Ա86���q��+1���CY"}޿~�6eŐ-U��}[ۍBY��f��Ku�� "0�����g�}V��/% �1�9%>'��U5$��7c`zb!��A��VcM����%�>5o��� h��i�#YͲ��Zӱ:::���g;6���zx"��`:�:�8�q� �1���@�&B!����Tz�2�U1*'��7c�2��şB�RZ�u��y�z��1��[1�1���[�S�V�i�©Ma���#���Q�Z7D��j�E�����:��4C��X,}�$Fw'+6J��i�l!�)$奕fl��Ɓ�X�kݼN�ky�Mb�Ї_T<�ō �2  c�<J�fX��H�.�Tҧ��Y��-�z�������^��QP]�7���R��?��n0u���P�d����:�L:�Z�<�p纚s�0ʬ)<^W�(�_^K�u�;Y}��hW�F�w5W�����?6�u
���C��ҍ���?���	m��������y5���_�sO�ŝÿ����GHgX��Ɏ�	$P����k ����ݪX�:�ũ���fJT��2��h��y�Ӭ�{q��*�.�a��1Fq
��6@74�ܬj<5^HW���ڝ$)�u��������;ɘhZ��Ŵ�Α��y�پZ>YG[�,pY��a��Lu�� d�>j}^�K��h3
c�#�Xi��_��[��,�D�AQcnoo�x��0��5a�B�V�kM����S��%!Eޫz�R���of!V�㸜!<4��L}�"�cr�e3����A@[��Ҳȏ-(�hh<��%_i<~��W��2�f�t0��o�),���&�����j����9X�`�ke&р9���2�E����$�\ˢ����
{Q"���<0��礠�O��&^���4�I>�]�3�In�]�C(����!���ݿ�,���wbb�<�8����K�l��ZR4Y]Fޛ��y�ߋ_�����|9�����~ܢ�����:7�t��� I�-ʛ��G���Y�e�+�и������bhd FFsu>Y���t�0}f5v�6b}i)�E^\\�:;�@@�eJ�[h7�u�d��z�rV�jo MM߄aN�	�.r[���F�#?�)�ѱ��fq��$�6���a���'�DӦUk���Da�kN
���-.8�;�u�j�>S���$�W�+S��2����4���=�w	�(8_·�'Ȭ&ʖ`�R?�F���=�qGgJ�%�!�Z�������9�i]��Lܔ��hfK�f�ЮB�[X$y��H'��]^X���լ���n-?�A���;Z��'x�,'��0b˟��B#:����=Ʈߩ�/B����|���Jļ�n�,�n�~t3v�*�?:��-�����_�-��������U��M��9L$����w��ى|���0���Ž[3�<�;ލ��嘛�i\'3c��ӷ�㤩�ݏt���8~�/*m&F&�u��~�`�d�q5���u.�=��b8�]�0��GP��dN'��I�$��q��+j��b�T��^��Mx��
�ld)�z���!OK�m9.~3	N��׋�-���|����A����8���w���+�T��Q�pRN��/PPҿ�=��
�BQ�m�3j�0�ex�	c�y|na��߾3���=-�V6���g��)cfp �p�l� �4�s�v7"7�5�_��6ӗ4�N~��'kI�%���kYF��3�j���MUr��M��g(��?�Z���3�a���IO�'$9�<[&���ɼ"C�.��^>K�[|S��s&��q)�h:��DZ&��u�vf�\\�ڛ(E����
�kd�@�*� }����'�Ƀ-�-���b{�[stv�Do�Gܶ� K~�s_[�%Zwn$�C-%<2b���P��db���i-�y5L^��:�h}s=S�v�|���oa�S#����ʄJJU�V��76c`�>�oc��s��LG��s�N�Gi�bw8B?+����5T�h���,���e��,am8�AkM���z0�k!X+-WS�UwT��r`	i鹾�t�)2��dz:�Vɤi��oe-O�-a�Q'C���$��b���������}Ԋ���>^�p��R�˞րF��B)�8N��Z�q����)|	5�"2mI�-		)T($-�Q���s��߅��7�h�����f�N5ʷ��}ve1Y�㜨��W��*,�K�H�wj(�na��z���N�UZ�+G�ɗާH#�J��������{�|��E{K5���T_}��j��4�>��k���{��q��t\��N�.��Ό��6x	�ͻ���B����\�,g��:���$�����:���Դ�ƺ���n$� �����40�� ����?��W�0 ��"��9qt��U+�1:�S����`��lVQ#�15v7n|x=�ƅm�HU�Q�[��ɄE�+$Ŧ�GI\?�CC;��\���#����i!�m
@`���x���7�9��FpB3�����r��>���	���i)վ����/����k0��e�NU���K$�Ȉ2�̗��%�Bv�M��"3�QR�^F.I�E�((&XJ6�Wf��t�qY�Ѣ&P ��+
��>%���E�w�6���EP���f<BH�H��e�� � �p=��d4־�k�ͥ<�9S���N��m�P�����/! !@޿��vn�_^�vi�'mE\�<}�W��~�b�V�ǝk������Ɲ���͸���Yo��(!�	�s\�K��z���F��̕�"��n����0l�t��W�daښ��>��o���'�B#lG����cH3�
��Ed ���jAW�<�5�EkwKf�Oݟ��;3t02\��ė=mY����A(�۫�d+K�1��Nl�,&�nWUbf�鉶�Q���3�կ�gN0���-5���H�qs�@�u̡0��y�^&�b�	�Z�]|�=!a(�u8J,v�\���e�� (�d �Ŀ�f-��	��� 	Ex�k6~��&���0��䱧��U���'!���W�w�!�,k��7��e�У0���!}�w�E�k1��rI"ۖ�U��W��a�罶�m�9�t<2����Km.��V\'�|eW�
N��e��G!5{ނ����@�K��2�OE�����l��b�ȏ�k���?�w-mɲ���(�5�܃�"��߼�|�YX���O��r������U╗Ϧ�_Z<��>X�{�*��؂_ Y�ޮ�64�!������~p'eb�� �ñg�e�{#����ډPP6�/aqQ �-�\U�����M��:��u�=2��mN�2V�l�S ]3�3@r�bjr<�&�} N.�2!����[�5��֢�������:fBWG+B�z�[>�z:cm�Yh���矏�~�8y���ט�" �/-���s0�8���̩e�gж̣&,[h��MS��l7|���Y�@���rKc����\Ӳ�	K���=�:foi��p�U�@��ۊIZu!�LdS����p@-����	_��(
���Z���2�"�i�]z��hf��`d�O!Dh�!���^�CHjv���63į�*�$7{�M��y9�h2�Y�M��)��V�{��"��*�@��x|���9��Ҿ<t���Z'�]��s˼��:��ۯǇ�>�ɉ��s{.�.�fi^+JxhQj*��i���VË�Y6a%@EyW��G�P{t���O�4N�4�!@��l�ϩ�;�G}W�Dc���93�L����ҚK�.��y��n����A�ʻaS�n�ψ����$je�Wt ���
!L�r"%�;�=OL+"�y�I{ow�7U��}X��|֏����`��#�uRJ(<��?y<�^8]@�}��*C�hG��9F-Z��Q7�N����-��Bè�/ӷ������jaQ�����'a�FEK6�&\�,-?33�Ș�O$s�a��O��d�fʣS�F0��+�
�B�db�Sx-�&�� ��~�g���>#�*!��4r-+23�J�o截p2�/�?�&�
�}P0���9�d��F ���7���
��Is�V�#Xek�
��xt;�!��o}\��`����$�/������O�n�K|~����Z��lุd����y�G�)U$����C�F��DM��ߟJD_{c���V�EooO��m��C��X�������%�뙸��s
R�΢���FH�N�Xs��K)d�x�r̴����ũ��{l -?�@���i1���a�)�IG�k�����-.�F���8v��7s�z����x�������q�����?V7!js4W�9N��=�fi��b��ז�폐O�Y&�,8��r7���L$�`���Vc�r�e���Z���V@6>"�"tVs�,,4����Tޯ�,�����70�L���l���v����et�K���d,Ɨ��+t�[n�^��m�Z�l�6}��ZZ9��w���r�Z0�am߱=K(��h�2�آ0�,����M-v
/�+�T�:�y�l|��,�. �+�)8L��#�(B��Cq��>9ƣ�*�wn=�9��s�<�� ��ț��8s�%��[���}#'�'��+�/ǩ����G/�_~��9���~��v���������2��PFNS1�����.�V�������G�^~mvj9��ގdVϤjom�4e0N~bL����?u�ǘ�hBӪ��I��H���[�����7�K����S��S�Ntz{1Ξh�Ǯ�ݛ�q���^��>rl(N�B�*B�\��V��r��+~E���
����2���#��O�z��GkC
��f���J�}Ge��L�*�;#�iu��Ad��|D����.B.a���D�oJ�*��2���uN�L�����	�O�%cJ�L�zh)�7E��Saߦ�	Se�\�y(�jq�Z-��ըE2	:Y�K&�__%��|z���p�~I��
wQ$�[67%)S���KZH����(��<�Fҁ�:��ڕ�n�E��cd�u��[�j���g���'��gOD?֩��O=�d�;w*�z��=@��>Eq�C�|�ͣBQ��܊ ��kx~�����G�Êe{�|:4W9dRd��}7��0F��:�����Z�i}E-���*B&�� ��$����ndΣ�%�R(�.L �����Z�:|��qX7o�����r���h��=��N"W�"(Lx��������ʒ��M��gd�Yz[XȽZ��������z�/���\G�8���z������d$%�(��H��e��.��@18��8X�T���O��3���>�
I�I�B�2�.�1K
A�.�ge�"	���A$i��ɵ���*�M��FjY��w���n�Ia�3�����;N#�G2)4�"���݊��2Rjif�XP�P�t���<*��:��������-k�0��MF���0ZH޾���h�g��42��r,<�p7FG;�䩞���s:3�|~�u�M�_Xc}[��A��:^(-�z׹p8�{��<s�'�G?.V������y�SC+�9��keq��`����h�,1�xSӻ�e���f��k"H��0��}H�>9�t�[!�S�j��m�3��h�]�I{�b>�K�̼�1����B��0� ��6��FcK�[���tQ�m�\i�k�����j�H��f[�xN��&R0�]x䡀�ō��L�[J��ۻ�X'���<�^��D?�e��A���(�nC�2�4�%S�}�B�9IYD��]H-/d��:L�)��պk��5���碭,�/k`�2���~�°0M��C��γ�A>�B=u.`�����O!�o}�=��iS���2��Q�U��E�*1��V����3���q��(0V+*ZP��{��*]fdHE_������W��g�l�ZY5���Hi�
����4���%J3�W�xV��?�wn`�ꚹ�ү #�Z����j;n�����pӠ��3<�JV���_�F��_�j����q�� )>M:z��Ɯ<�/VæC�K���N�D&a��h\�V�P���&Q�����s)����+�FjoZQ1��j�-�jrS�7k�ip�Cs<3̈́��I}���ϴ����к����}�ٶ�@�M�bqq17���k���,j�,��� �L�
��%�����)�׺����¤l���KF �]k��`�Vn��F%�����iM`~�M�z*4�g>|�wc��&�&�sn���}h�B��d�S�
X0�ݤZ��"b�5�X0UA��a,�ʚ6����>�<��i�S��R
�˜�z�S<8"�sܾ�&yb�@�~����?�|?Ү��ہ��E�����7���}}��ݗ��D������ҤX3�)q��3����ή��ɻq�۱�bd��0��;��&�y2�����'v6�oʈ;S����R����鋳�⥗.��]�<2�<��F�X}�?k��s�-��G�
�m�qj5��:<؊�g�r�6e�N�p�	(Q���Z�l����o�&��_Ilg)����V�uj+�������R1����_�M���-N�����\��U�G���bRj��[E�D�ݵ�F�u�u�(��+*[�@[�~�{	��ܷ�Q t�:��Ʀ�4��XAK�O�Л�ad��O��@�G� �c&Π̳�i����;�Pb�OB`�.��<�6��9�\��>��9��٘Y�	�a�x{�6�^CH�66r��$`K��~T�2��Y�]����X^ZN��֒m�n���,�7Eø�����x̵T���2C%e?UjB�\dW�B�������P��|��s/,�u�f�X+���A4э���;!:���cE������Û��۟Ʒ������XXY�'����Q8�%=L�Mh[���f��5;	#��:|�MnU %��	q��1�Ԇi9��P�%�:�٢=�`d��=^-0�b+F�Z���^�{+K��υ�h]ϨaZ��6��:	���ؿ�Y��-Ph��^������9�!k�w�a<Cʵ,�*��dNh��4ұ5��jS��"l	��g���}+~���d�� G�@E���*�1���Z����0x#c)p�ׁOno�LY��+PŪ(�)�0��U����b�sΡ4�>�'��9������z}nӧL���Cɪ�x��baD��?i���M.���)�hy6���5�'��mjS�½)e�M��8B#�'����8������=�&����q�XS�5
k�߱��%�{:�#[p��ٔ�s>��ZH���ڕ��8uf !�Gal�d���639�=l�����j"�`�.�K�݈�isrf>�[�Q�~� c����$�t�=>��Z��ֵ����J�gm��@���jB�	`�a������b�M�/F-�Vs@�'c������ތ�%����0}��q��pt���냀��*55�X-�&Lc�Z��}w�����t\��f|����ug�϶���,�\q=}fƅ�ZD'����ѷ:�d�l[�Z�WC^�LmCƲ
�tK��]�N!D5�7��m�jZ��B��O���T_�����@��ɸ��H;>�v�Z�L�K��{�����X�$w�sSf%<��L$S!�/�%���e'8L��õ"
��+ŤQ���u>�v�����䧝O��P�weY=� J���>�0SF^�a]=�ٗ��}�~,�����JVKV0r(��.uǕ+#y�m�`|Q�ձ�Ʀ�����||�޵x�����:��/��/@|�V��^�6,��'����m��zƱ��!c'���ҕ�����+�|t7;12�ˀ������`@8ȃ;Z�����0�t&�J�u ��^��V��j~��{��*Ү=8s�T�95-2���� >΃����a7brq�p�t�5�Dw{g?}"���W���,�D>04�� ���9o9�rsgh��~t+���?�����A��w��H\z�X������j�`�1YV�jx�i=l[�Z�hZ@����j4�p����H�6x��桀�.�[���j.��ZP� ��Ң�v�����

�B�=�����v�.k�����2�V?�w
�Un	��*�-�D&�9��	��g	v���]�� tƶd$-��~:��2E���f �w@9��H�����K��A*�ʶ���`{޷c�yER^�3��f��R�Yk��b�=��k`��|��q㓛1�`,�d=H�j;���{j�~���v}���B�M�G^+T�"���i�x�z�@74i�)�p�E.ʰt�kp��Ώ��*�ft��Đ�y�+YQ���#��\�x�9�[���ݚ�)�<Ւ\��� ����ͱ�_Z��fH���%�?C�m�'�8iF[@����V�w*�=���7'��gc�ɭ��[ٍ���X�����a{�H뛲����'�+Si������&�� Ak�`��������?����X�����A}���>&-*#0��T�\c�B1�
Q� bZ��Ⳙ%����j��j6�����a��F�� Ж� -�E6���25f=��(�h��`.Z7V�"�\��.
���Gu"Dkn��ZC2�A�ҟ��X�`�3���?�=G�˾dp�U9ʖ��\Z[ڍ���Jk�\��ᘵ�
V"��-+`�!�}Qȥ��F7a[X	�ƦG'�����Ų �ȘT"˫�q��J|pm1>��K�����T��XK�,hǘ�偍�\�� L�	�9�}���A��N '()��Ҏ���a�f���Ps��ז�טö�Jp�X���i�W6�(�Q���s��	�(��tM���	�?7
���a:��$�`�F~on���J�4�EK�[�ˉU�`}��`:��QA��;���H2n�{腻\�Z���OZ��}����S�&��`��/yF�苫O��o.�"L03�5L6�(<|���Xd��@d���52fr	�g��v�p~³�|
�yn
��4�Hs��×�!��Y����ũ�J�U��M�u!�g�/Z�Z͟KZ��;���aS@#��V��f�َ�$d��*�J&#̻��=Zi3l��i�T^k�ʱ+lj{"�#m)@&�Hв@$�J&�g$��� a��+�����o�]�wo�6=�`�W,�-1z�m@�X��li�K��]wUvF	�.�6'\	c�,,e��"�";�'r�}W�<g͚�k�e�����wtt@o��|2O`Ա^���9��bY\M��f���O\�Xyb"R��l���"�¿�ccu/NƉ3���k��ʴ��{�՗��K_�������a,j��z {��HX8S�R�T L8���prM��`�;�ß
!��[��N��j��}s)���Ape$�ӬOC�l�]U,�	t)��2x�b�x)�*-	>�[����E��,�	Ӵ*B�������e`�m��QR���~�m`_�Ɨ�V�N�O�E9-���^��F�����Ev���m�fV8�$��j%˺U�x)
R�%i���e�>6-+�${o�;ф���Z�\X������*Ε�7i$]H�V�5�8�J۟��k���%-�tQ@�ӝ��d��VZs-��pGtY*-�ql�1zz�o�3�y���;_�R���S�ܳ�gMOi���'=�L�-�E����M�r�6�^*��O�I�-,�¨�'�[@]�/�L�|�����
�v6.�d$�JH}a�!�ףb�h�"�#�i� hj�j����+��/���˯ĳ�<� ~��+qr�3Wb�XC�;��?�����*'q?7��������p;���vEߠ�/��TӮ�x�g�����t���d(�յX����S�>���ܝ����8�+��.��cg�"�����L�����S���+I����F�0a���\#�6�c�4r]���W����=i�
��>�gF��2�!��x�
�C�]>�\�w{��U��K�2��c��B�؄E��Q *�Jn���3	S�X`��,t�R�c��( �Is
�L��0Z����屆�o���Γ��ߥ�Gnq��Ϡw�o���z�ss�V��}�_m�N|��'�����K/?#C��\鋋/��`_Ω%�����?�~;O*m��iO�������N���-���\`tcZ[i�Ba,�1�վyƙ4��	4|�D����7xp.�ukjU�r�%q���a0�o��w�2	�����NH�_�\<�����j�ގ��n��Z$;>�x.��!aX:��93�f����4��d��U�Ԏ	y�L�C;�\9-<˜�F��%\P�j\�3�OEwwm��%S�m�9�L�諾ړM� �e�>c�f%�d⺘�V��̐��B�$ |Y��}��z&��v&���p)P2�Q�\���S9�b�
\s�cn1a�ef�Qu�aK����wND�!�"H2���@4��[`dP�r<�L�ɥ��	_�Ґ����)L����ٮt�:ϲS��G��E5�7�*�,%��-�m�|�4��K�B�2ZL%�쿯�~�,� vT�>3��Ա�81����>����Ln���J��"3a~���e��6L��?�Ɨ��|tw��hbrɀ�*��4A�<�޴:-������T8�F.��¼v�C�#p�����V�rMm��1�od�+3Ã��2�D��7r�ڇG�~�k�ƩS=�`���Ec���k��	�Ԍ�w�r�Y�	�h[����"	!�$�)���簖/>�;�;���g`�M��8�$V�,āas3!V����S�"s��@߁���Ӏ����3�É.�n�W.d� �O�#�q�Hx��dP �u#��"����q� }3&�t@?ĉ���:5{�'�Z���3�E?G!�d-�N�g8޹4�Yh�0�v���[:K����f�\�L��9%�^�o_�����V+�P������v�x(`#�ZG�B!u�t+�Zi�km#;$��(T9�^k��[�M4!R�����7��8>��}�br�AB;�V3J��̺���� (A�[]���cij.z5�LT�hl����6�9����� ��<:ˢ��*3�s�Ͽ6;�����?��,��5Ü]1|�/Z�*�Ԋ?�u���\��D�a�Ņe��ynY��a ���c�zZۢ��-��g���eB�t�����a�9�?��q�8V�U21���8uz4�($���L2 װd\P�R[[˼�.l3��k���C'��*��W�ދq�l����R��P��6\p7��5�7r���b2�h��P)pNbB;&[��h�QU>�0K���i�(!�LH�m#K�qMf-p�ka�<SM��]jk��d&ڐ�p��{�Bhv����.���w.�r�t���*�dN���?��NB@�8a��{�:�8R��KZ@!�J�W?��ȽI+���K_]�X
-����յ�t��
� ��U$��F��b��u��9o�w�ֽ�m�{��~+���n��h�l�������9�C�tS�!Bɘ���w��������4���1�{w����q�:��5�]dE�����㌭D��w�6���������W��63mM�����{5q<������	�tS�����V_�N-�9��j|��	29y�V��n����D`��
�6 �����X]�+�������}��1�͕dV����@�;w<��,��o�HY]w�F�����I��ۀ �����q�cq��p���#�_Ţ!��2��	�d1��ɤ�gL�Y�h3���V��4sKY��9�M}�QGy�:"�f@�ԧB�AedS�2�E������)D%ZM���L��t8V���9*A�c�l'
AQ��S=12���Z_�]�E��S�r�GV�3Ɵ��7�G˃������ ���̒l���2H�r>M�O��5��ү,�>��%��a�����i?k����"�Bf����`nS�V3ژg�����x��c1z�;�x��m����=u�i �}�f����B^��
։9__^�*��
~���JLL��QN�gUZ�,-.fp���.�Z���,)�.mDY
3��6��gp�����5|��t��ޚ��[�q�;1��k�4���Cц�9�N�[-���U3�||�{� _�ue�b��[���9Q�r �ry��r�( ���b-�0I���c��.��~2�W����_:��B<~v ��0��亭�L��%��Ƀ� ��Z�,�
V��ig2�>g� ����И�`�v�&�8i��Jtgm�06����R,��6W�h�J�au
���k2�K[�8P�dl_.���B�E�O��o),\���逯Z��͝��X:���E#��D 
H�ʣ���h:�&i���qc."3*R�D
�̤�8b�"@�,:��ºН�C;Z+�_���Y�f孥�L!�@��[+��P���,�m�"I��s�S���y�|���wt�+�>�� x�1�?}O,�J��$v��2�a�$�j�j>�HA"B����0Ug_WT:qC�:�k�/N�=��!���х����)`�3��怋Y��*L�+��&Ǯ�6��
�[�_�- ��^�W7r���sZsN$S8�B8�f/V&5�~M�={*F�u3�h=&e"�/MF��B�-N������ϦbzE�N���ȡ��8{n4O�Q��a@�>O���< �Eu���y�4>�3&��x>�,{��@յ�Z�(��\������/�\ZJ����Mz��g93&E��-2\#�g�Y8�QBⶫ�A-����I�^�s���,)�J�/��}�1m��c.�]��~'S�»P��2בg��V�Sl��%L+�<&�J�'}I�Ge��矟�{�����'_1���«��a�$҅����c�D��/,rۧB7-\i�du�>��2��Riܾ}?�m�����,���co3�x�s,�e�������6�c�͟��}����)�u	U�c��uUX���mo�����aP`&k�Z}t�ͪ�._$�@��ߪ_�����Gws���#]sۉU�`�����y��	U ��%��⪔�������E_���#d1��>zm<r�R�?7�D�@�>�ccm?p\��n�o�Ɓ�X����>�h���_�����*ת�u*KXm����c�+�Z��9�����%�=�(5-��:�f�Cw˄)�j#&��&&L�z�,���+'E?Fk��<kU2�o�p�f�s�Br@�^jokG��3�j�OFSx����M���H�\�3-�}��
�}s��{�1�mE �?�状���c���Ei�����V���^�5Jx�����*�E�G�c�f����p�M�΀�G�T���Z��h=�!�Ȁ�h��L�RP	�շ$����m���o� >�v3�_��se��	�������㹧Gi�h�?}s2f�i�a����;17�q}�~�TȌ�Y/�P��-�;���2µ�`'�����,z�o]J�믫��P�&Y0ߏ^�����D;>��,�&A��+���2�B
m�`ii)s�Z��\P�:1GA����6��ccq���t&o\����b~u7�������Q��\�%j�'G���y;iN(��a
�.��U�Zա5�^���XIP��������5�r�����7�����f��ʠ<K����f �T����TN�^B���«e�N^���jp��	M�(��)B!��cw>#b
���=}P���_�fthA���S��42���k���#,{�Rhh@ڗ��IuϿ���W���}�"56j̀w|c���4.��/��~x�(ĝ�i%�7�atڲ^c�քQg?}i%���O����H� l��>��/����g[���M���(��hj�U�Q���7x��u�ȓo�B��{⩁4k�l��O�``C��YڍX߄��{�y���%�{"�+�>����2DĒUp>�N}k�W�$֫w[�ĵ�c.6>$�pL&����mh��Fh �$���J%N��d��������������Ry��0d?OE���U�k=p�g~��Ź3�3���B^8��H�wT4�5#3�kB9X�����twr��]],m��n����wSr�a*pCB<�*�`@X��ڞ[<�I\��J��>�	�I]�V �$M�l��:�/���`��Z��P��#�p��LJr�E�5'�Rh˽��,�������G�T����Y�z#�iᡧB��HE"c�SE��G�I�Y�ysk5��(9)��@-
���[�@����kz��'M���пV��x���W�dQ�}H'H�,�7
���x>�|,��6�4u�%遫��S���8Ċ�	H����P�F�U:��W��B�z�to_O,�-���3����{!�V
5#`Ҝ������Ņ��
��ҕ˯�af�Ԏ�����,���oh��a���Bq���hi����FMf��L���N�Vb�DٖL.��=-�����'�Ѿ���k_��>�7�ݏ�m1>�FΝ?��mq��p�&��;#wL��ɜK�-m�-�υ����/׋���R�L�}M��@䎨�P)(N
�k葳��IL�y�OA�(�ơ6���1�w��ZX�(�Z$���8Y6���k�點�"�0C��(mɶD �G�)��v������pw3�e����˟�~�����/�Կ!R�=�%�=7��"�F��2��粴�B;�˱AKO�-���*��G�C(T%�x_��/#���(�J�+(9����MӪ�Uc(_�U@�f�)#����q��%6��-$���{��Mu�c�ܮ������7����_��_~!^��s��ի��>��h���,(/ !5Zy����"s-��P)�+Ȱ�!�S&*8����j<\^�~�.5W}���5�����6P���T�r��0j9!M�a�Dȵ�fB,�9�}��;`Q��X�[K�[4P[|����;�/>%�yƼ�+ql�z3F ��Ѷx��1���A&� m�81#�}X�F���C����)eT�2F�Tq0�ap'J-l6��a�&'J�Òh��@D�ie�����%5�������k�m��0L��6.�&x�Yimx��c_�Y	PxO�E��g�	}�o����h�Tf�����c��lO��&���~)Pkh�����F;���edp�K�x��	�T*����y��@����Ԛ���'}e:��*yH�Ah��L��տ@+>�>+\GJA%#ԓό�9��_e�M�^�� d~�j.�ܤ@��kv��v6����+�W�ĉc�P��q������*6D;�mh��[���Z*�7B����.��6���uE�>w�/^z��h�~��v��@a����O�!�����ZМEc�qv�bk�� L��Y*���!}��ۈZ�5�3!D7c�����3�k���o�g"� d�����L���Ocf�s����`��<J5���|���0��X�+`R�a�{����F+#P�\&��N_K���W��4Z�z� �2���7mh04_[�������|8?=�>C�ܫC^�32؁�h�6���Hb�4a!��PA�Yͨ��U���r	%�'�ʀG�^�����B.��yZ޴tE�'m�����������K ��{HD%��XQɷ�[�[�8j���kڡE%�cR���\t7e�9�+-�����f+�w�M�P�������\�۹��ԕ��X�l�UASAH��0D(*�=ޮW�E��Z;��H%����`Ct� 6���{1;����N�iג.����D��"��A��j(��f4�� L��|�T�>},��H&�+�ilPDe^j�����&JP3ik5��S��O�ύ0����G2QRC߉yKl�A�����I�^��F�����NJa,��啵��ߌ�����]�C����Q��Y��.�"$�xHp5#JX�&e�An0p�
��-ӧ���� 2�?����	���n�/��l���2��s��Eț/S3��H��{X�%��j�?oV��u��2�o���j�z���(,-tK�Il϶�3d*�>�����i�L8ΰzZ{��n�0��n�꣆��f�}�p�7��4�\,��Q��f:��W�U��iٹ����V��>BX�ؚ��{-�~�sѢp=T�V�W�������zH��C������ d�D N��p�����և��s(<�6���Zv!���j^/oi(���?l���!Pڕ+'�ң'��%#��凂/�p:4�u�DX�.D+�
Z5�3�[M6<|2������~�����ĥ��P��^:⦿ �Z�����ݺww6�ް�g��3���9�h�4�
�Ȁ�4�"�џ�������{��Objj:��\a_����};�Y�D�ot΍w�q"�������)���X3uG�ސ5��l/,.�Ҳ�-���oe��k����� �al���En
cK[ ��_�JG�u��{��D�`���MF���q7�;�մZF>KΝV�{����s������;��LC���5п�e��gBi�m�Q	�y��mƚ��epY�W��Nj/E3r�!m�T~���W&(�t4�Z��1�w�������I��ۥ��
�$f�,=?�U����Ĳ-�(�!����n���bT7�Dk�.��Ra�>�R�<$R�~*4~&�/;%�A��X_]���t9�ѝ2)Xw�
U�������������l��v!�(��Q[��ã���`&�>�k�o�u���U4W:`�>O���",i6j�ξn �iHNn]45tǯ���ů�ҋQ���يO>�(��0^}�B��k�����>Z�U�����}>N��|����V�ψ�A`�Ԫt>�uL�L"�l�h!Z��sd<'ԉ��e2]�uS��M�Y��I���_/��������cS��蓖�l��A�E3��k�^_��[E&އ3� � ��=᜵��^��wB���	����JS�#��'�� ȃ	��-e�q�g۩Y�6��f��P�~po.?@;�]/%�C���e;�i�D!KK��{�fX��XB	�@ӇL���p��﫜zR��$�/��[�Z+�Z�̹�e;*~I��� �ҷ;7��O��[11�R�o���UЭ�q'�ſx9�\:�����g�J������F3ض\v���߉����oca}wAEW�dV��������E+��5V����`���J���ՌF�֧��?D����Lި�����ñ{�14Ԇ�f�/���ֵƕG.�sO�
J،����G���9��եXXX��\a�ar,���M��\+��<��Jo�������o��@����ɛ�X�� �D��L�����o�B+�`Y�$�����x打��?��h1��dJɏ�p?�X?K�碨�!�trd*��,N��
C�M2��S!�y�L�����H9�4�3m̖/M��+ia�[�N�@ߒYy\P�R�dS��	�S��G��e ����?�4��ugZ��R�-����*^��*��B��ل��ki����L����E�l��}�}�� v����Mje����ܗK�Nf.�}�?�}x}���,��Z1�U.9\�ӝgQ��Y�u{*��z��* cӠ����uU���7_�/��x���O�œ/������<�]����?�����_��⽨n�)ZG�%�<�ow{#ݍJ{+��k�+��d�+����e*���.��Z�ޭ��kկ��o޻9�����"&n�&���ƒ���3g�x�^-�����x��[�RѮ��,�555������a���s�n}y��'~�w�A|�k�F���[[+�q�1A發�������*,6�v�����'��o��`%���������XZ¥�e�,�CJL���d�AP�n.��S�U0�f$�j8<��8x>7Z�Ҿ���jd�l���̘	��p0�Ֆ�m�4%cd���{.��/yT����0�d@��~i��~'<���ޔ �+ê��}ꦀ�h��$��~���
G6Ry��N�0R���
5S�2-���>��`��"��:{����z*������06���˵
�s丅�Xm�ʽ���7��RI��e�-��Ew����x(�*Ii�h���~���9>~�N\�v#�f�3.�\�������կ>�K[���jl�v��2
��.��c�*�����G��X�^��fx���9�BocJ�����w'����F�$�1x�h��ʗ�� �w'@|X�_��_;���D�vFO`��f$څg��
h3&L��б7UƊA�[{����z75�FkGK�w7���f�.�ä-��SO��3�h��\pſ�ڎO�{;�v���*�9�T{WW���S�ֺ��_|'�=���La�u���1t�6Z�HGՒ��A�����s=�KO�̭3�M�;��ik}+&�Nƃ;��a���2d�QAa 7��T��á���d���7b5a
-���fK��S �1�e2����-"Fq���;�sF-�caf&��r���E��dĨ��T��'%"2^�/#q��ϽF�Ѕ��֖���a�]��>�o�Up�>�����F���DkNh]�����Yޚ��?N��zY��.}��\���54�Vk�>�}�I*F�p�,�K�� �ų�R[SK�?:^x��ܵq��b���)>�l�0�����ʫg���dJ�Ĥ���`��2GThc��9�7���׫�.?Yra+:ݑ���%(Z��a~����4}O��K9���{q����cq��o��_9����1N�v�B���vL���(�̨�������mvsQ�C��k�c�o�hM�eԥo�#�)�Z��J�-�GDik������������t �z���Jܿ� ���b±�\/��jV��[a?��h��s¶X~��k @�sݭӣz�Zo�݋������?��3Yӂ�#����ݤ�X���ej3-�L]\��:��%��>�;�����#�h.����-PHU��d�z�-P�!�W��D���q�C���	@�`&Ӎp	�hO��n�����tZ�:�+����6��~ J�H�	�|U�~J���z������mB�v��C=@i��7�Q�[y0�c/5>k2�W��i����TT
-c2+ƃe^�f��yu�����`\�x>�A�}s*����2��d}h��<7�i5�AUs��1� �|L�P`�����#f����y�>!j�g#�5Yè�¥k��r�>-;m�X��bzb�~�0o�����M�L'oh�����"�\T9�:Q�ʷ����ۈU�X�z��Z:�$�#Xg��sվs���bv|>�it�Lu��"�ƕg�Ž�7cc�=8��L���1�:�Y��k��X�G�w'�͏ޡ�eTM_`�_���������wbRK	��xʻ`�r��
�P	�%�BE�(���P�ka*�Y��s�̉��4I߀u
��́���Eb��я�� f��y��|��:~ƸC��aD�� �0�T$5��sqaA
�4H��������Ae�Z����mdX۾
��h��li��-��{�N?L�&2|_h�:Zms=¦�a�T����� ��X�L��[*"O�A謀���qN�ؿ�[�ܹ��?�m��ȝ�KS���[�J�3s	ێ_Ν��g�A��4_�ڝ�W��*a�0��9�=��[̌$�gi8�z/hO��DcCs�[�h�ᆆ���*r���)w��x�)7^2�����\]��E7cee�a.�SHcZ�&��
�S^���T� ���>�\�܅��C��;�r�wmt���>�dL�K�����]�h_'��g`B"ɤj`̶�l*�L���|�k@���w2���j�7eٻC#Z���lQ���3�Hɓ8���V���jV��M�QN L#�c�!�����	Dn�:��[�0��<Z'����ku��2���⮇9����?ԜB� i}(�2��yP\\hDPkj��B{݌�����:
���4#���:�D�R ��J�NN15��S�o����ہ�V$k����¨R�|�O:�9�~c�ވ�)m�XZ�_��K�����U��v
�ǽl��W�rEI/��82��Հ.F(�?s���P�FbU���<����c���y�t����<��A����D�\?y�n��
�tC�݉ �@�@��o�����UvQ���H�W�5Ji���sν�0�s�
�tfj%y�A�2Y{Nx��9`3�w �(4[W��,.�fH��t�r��8��v	Z4�N/>�~]tŕ�g���;��<�Ox��%tB7�B1���0��h_�q:̛iI2��8T�Cu�tC}��0h�p��cv�sq�l�uKY�H��5U�xjJ3S�_"u�[Rv3^\ண?&R�p}>[Sn6��0�4��<_����<�x����ne�c�0sA��$i��M�ѵ	0����c��`�"�z�m��`���-��˵�**h�x�s�����B5o��f�-ڃAJ���50�t��i�#� ���*S49���5m��$i��>���S����j��Y�C�.�V�4sQ*��,���.Z8�RIz���X//R�ο�^+��*K�#�S)u�zx����>�Z��],k���
��AcJ�;4tE�j����
�VWE��Z>��e����]{���҅��t]~�W��O�s ����֟��*�f�*P��R�+�Z;y߁�-̢'�?���'ӛ��Y�t;�Ź��_�'.?��_���w���{&bp
��&^VS��*�|��U���7��+y⡖,�������������i�m
̅#�Č�q��'w������[_��	p>�e��ds�k�?�ٍx���o�b��/|�R�5��l`	�������x��g�Pً�~�R73a@
4��8�I�7?��ډ�=l�ֺ���W�GG��K�P�0����u���m�0��0��c��KH�	��˴���q��l��g��W��~<��P����V�����ٽ�~�x�)�.�W�c�DwW�(dt�v��n�Ǎ�������G���\G�1�MO3A��]�0��ӿ:ڭ��[a��������eL��ؔ���� ���l8_�UY�t�P0�.��B���]���5FH39>�o��`4��'�}
<gl7�i�#�z����X���{fP!��[��B�F�mJ� 8��l ݋���Ѻk����\z��k�)��52�m���=��M&(�D�:0a����
/3��]) SV�w�_��	�B��,Ս�=��.��۟\����t��  �G�"tβ�Ȗ&P�8A�0�q�(����s�kErcP8ϝꉿ�G���.x���X�޾���!��{߿F;Mq�Dw��o��������;�^B�7s_��aMZ����;�����8�����O?s>{�b&�^�hZ�Z��_�o~+.��. u-0���=u)�>�|?{�&}���p%����?���ၮ���������cэ���a���/����|5�}�\���V�E��{�b<�"�r���w�k�⑋��_��W��_x4.��!��y�ɳ���w���o܄�����������_>W/���޸x�'>�ʕx���i�>�t�5�����g���\�'��'�����x���KW��}��\�U�����F|����3�㱋}�3��|!^���hm���Xl{�&5�@��c�M%+��<P�	f]���y���@	���M����xnG1�|jr�ܔ�f�)cR��Җ��-reh�]����� �XĎ��q��YAn�}i	�]"@��YxV��:H�!�.8ª��t�B\~�L���#�e��J�=z{h�=����n*a��zJ]^�D�p���Ņ�e���2�����S{�_�~��E�ܒ^��Q�l��`��jY=�H���M��5��w1+Am���<�?������N�9�7߰l���Z�}'����`�6>|2���n�_�ǩ��?�?����\G���_χ~����w��~���4��>�7~x#�u��bx�SA�<���g��������a���?��-hZ��:h[���orl!��Oߏ���|���~;��ں�����쇌�6�����ǿ�V���v��͵?���F+
3�5���т�\E���������7���?��g(40߻IW0��R�������f�?�ߧo�;?��|�n��j�@����B?�7n�ҏ����Ż �Zx����u�M]�ʮ5���w����˿�et7:�ڣ�":r$s��#:*p�$٪�-�S�	S���C�}]���Ҳ��)}sx�yl��
�=���EnsKs&|�(�����M����F+����Gc������c����bh�ٱB4O�pe
{����_�����	��k�L���HuSXε���L�����,c�i���X�6��isGgg�<)��(3(����ۻ����S131k���tC�.fwY!K��0��f������ڤ��lTS����хskMs���k<&�G?�7ƫcز�� <܍���x��O�g�:�k����7�cj�!��Y[{`�vB�w߹�?[��c-�1��?��͸q��׵�5���:��.�~�f||m�ɣ��W������w�O�ۢ-�vݵ�����ѻ��}{�hq=?������+����;�u'F��^�7^����n�������x?~��b,���R��=ևb�?��Q�C]q���x�����{q��jL����~�@ӱ����w�C1�tOK\:7�y?�������NĹH6�a榸~}6��@+�_�^�?v2>`����⃛(պ�į��i�����&��4��/�t����Ν�=15{Sq��P�ۇ������()L����J�7o��pPR�,��ZCݙ����ϴ��eŀJ�-P���Z֞1��S��^�
����³�=142�����n�u��n���|_��Yܠ�X^XF�5.U��͸]k��Ok$���s�MO-&��Js�8gq���/S�yv�w�9V��ι{zr���0�0*Q�Zk[���H�-Ko�g���������-gɒ(+P�"9�	䤞�����P�*2�~��op���(���=���9��s�\%a�Fug֬g�GX=dI1tB,�s7xp���4�%�t>���P��TZ�ӿk1nGgR�}��2�}:]��)"�!�ho���ee9F�:�o�tTDm��~��4[K{ʺ�:����:ۚ}�YG[�Yv6#�C�ll�0vZ(�be�VIX���vk#6<�h�C����kU:��jR�V�֊%}yLE(f�uq��]L�ԈZ)�k��^��-�j׻Yצ�!�bq�,n�ݛ��3,��/��ne�ϥ$Y8��b�����]�2b�r�z���eVe��-VM[}"i��^Y��]�t߳m���0yC����Ү�NѰ�jB�O��Է�~��n�bPS���j�68�a�+r�wկꐔW��$����#ʻa�;�,a�X�o���[�΍كт ݬݽ7X�2�I�}x=k��5VV�)�u��Y)�����M��m{�Qo��dQ�Z�D�*��ƨ�M���y`����|v�"Ѱ��-�T �n��7Q�`�R��;��Tf9�,��Z�V�]U����:KKi�}ayU|.WDЅ�+�ܼ��Y�&��>��[�Qn��,6W�6/�`�?Y[\ȸK�5�p_1���l��A�J��.��"ޙ�%�Ԯ.<;C��dw6%0u�O0dcM������*Y��,K�ݻ6l�d�?%�Dg�ښ���d�3�ᾛ[>i	����og��!,�EjM���u�i�Mae�>�i#"QD'��v �յ�X��h���/Oح�h4i?�J�_��
���;��-F��I]߳K?�m���#5v�ԓv\~�B�d���"�|�p�
֛������<~��lE�p&��߳��>$-�^�d�OZ_��b���#D^.��&���_��k��I+�:�� G�-r�q	���+˶��cO�w�{S�pC���g����˂j̘,g{[%���
E=�)A;���Oڑ'�LH6� ?�������%����}_t���W����O[EM�rEit�!�4��p����{v�NF�f�v+��s�I;�dJ�n]�����¾��w��{��mV\�[�>g=����:%>��*i�)S����1�eϺ:�lbtʡ!����B)q)�I�kl�m�������HD�>:Dl[!��}d���,����uMV��оS%���܇�A��#��Qʜ�=�Ҷ𖕄�J�&�i. �>���4e�ȺZ�G����8�`K�߉����*�������`��I��r���%A�9���ZV�@�ێ�< �"�'�$��}1 ��K�$|Pu��^��_�	_�b�"��$��*XdW�`&+KR��~R�nͅ��� �9%^q� ��FF	+�����b�N�������YgSJJ��uL����c	�
�t����;u����9)K����V��Ȓ�%���KJ[v�ĭ)��$&�A�|q*�h����C��!|__]g!��00�\d���ԗf�.�b���v$����z:D�Hܙd[cV#�����ԑ;|��ˏ�lN�ik�]���)PC��:��Bv�P����y��/�>�����#�������ѪS�Z�H�O<v�>���������;<�m�D�*�$Ȓ`3�h��:`O=q�>����'���'��U~L<W�j]	n�	�����A;~�G�;��aݝmB)B����	�	sbT�&�������>%(���x�z�Z�N�.g�j�΋D �Z�d�P�@t&�"#�R���+��n<-��īk��,��Hl w��~PN�W��a�����Γ�1*ni��u�k95���M-)ki!^�ނ�C�8�J�ǒ��oV���E	���I�[҃��]ؚ�Y�Yf��[��aNL*�|�� Sc��hY�Mɏ,� U���"Z�Q,�B`���JĐ<ɨ;�h7.����y,���Ⱥ��>w&?�������%��}li�R���쀢cj~(Z	? =��^�-��d�ˢj0Bb`��}�i�Dc��Yo;m�I�R,d��?�Z�/�C�'P2���p�Z��Y�����7D5���'AB�����~"��q��5�Ns��j�%��'�~�I�3�O0J��=��M�K�i|�Ԫ����@щX<$��܋��L�<��zq%݃X��%��Q��3�q	4����v��
�gl�@�l��Au/��h���65��@iZ'��q��A���,rH9�s�,@��/���r8��s����	��9�j���)�k�B{	��A�5��T��d����b�zC������$�kk�.�dwR~C[K�`_�577Y*��x"�F�(�aP�lzb�&
�i�S�dL�n",'A$��!��VO{��̏�|�켄��=^�I\�{�K��)-A$�Ox��JTzL�3˵,=an�Z��Y9$���?4�L4k�6����!YI B��at]ߓU l�ma�K��sg���9J+ �DYJ0A�<)[Xor�X,I�d�Q>�hئ|�=9�z�H��Jq�������n�ZnE�J!�D&�u�[E�4���H�vC����W�QCN�Vmi�}ۛdAv�^e~�`YQ�Ů2�B1�!��|�G��[�.�Jz>,)x���^.mm�
p��$`�;�:wV�yV�K�珈T�9#���mA���%��YY�|����</�@��qC)*櫈�U2;����e� (��ҸKis�,�`_Aн(���A1�m	Жe��W�ZY�Ij�X�~�c�h�	�D���Ak%HTZ��D3YS�,�e�X���d6|$~��� ;��G�}5��T������`!۞&����^CBj�剛��Jh{��uA�u�����O[V���,!�����%$ª��G��_��a�YҴ�i��P�A�:��05��c�_,�����y!18�1��KZ[mF�����aN���Ԝ��Y������ny�X϶C�C���̼�^Y_+ڃ�lZ�_�t���s]��{���Y1I�����qi���������G����!�p��ՏJ߁13��h�brt�n߸c��n�d�`�׳�3�Gfm)�s����Wo��]��w��K�
�D���ۃ�1�cH`C�G���}�nݼgc��m ������4odh�b&k���}�7lxtZ�@~ꪯ�]��ltx�2�y�:�s�>|�C�~�=|8"LS�VVr6��sϩ�i�����+��{��w߳{��jC�S��2�)��8�I����������ڻＧ6��e��~2e������]-(	jA�b�g�!5�1�g�@M��tX�1�袈uC	(�>������d)u�(��R.��/��]��Њ0�yx� ���,0|�
T�tt�{zAW)?W�_��/�]�>"��'�t����Z��镔Ɯ!��:s�L�+"8`�-��LMg<Do�|�ds�fV$��K�:G1ה�F�n��q=��m�KE_UJ@$��[�p��{�4�!�[-=��x�8�#̇ i�yL=���t�n4����[��ή�$?+����g#v��ӂ !i���5�ʔ�'�O� ?T;���j����DT��r~UV��v����:�6�}UU0C���%:����t��0uK�"!�Тk	��������܌�� ����ɢ�M���mm�hMA�\~Ŗ�����P �IQ�mV+F�+�����BJ@�3��lK��2�l�݇���D�٦OFO}3[�d�&�ԧ ����
*�|����2u���tqiN�莟X�GV]��,��#x)��׹%߉�l����o��Hڦ�s`�O�p�ڻ�~lqa�r++�D�
�ʯ�s�D���fY���L���!C��JHcĶ���t��Lɸrr%����b���5�w5l˧��c�㒍�/� P�Dz� X���YYS��K_����ۣ���n]�Ig�D����&1D�KyvaI��u	͎an�
s�+2��67��פ '��5=���z]�,ѹ2i�ߑ�ج:��]a
���-n�:S6�`\�h��S���y��n�ʤ�����(����W�]1H��zPWs���,� �ӳ�,|���&Y]�[���P@F�f�ڗL�di�VX*�VK5��mhD�B:P�ғ�7pб�d������d���B���0��'R��^Oy�ξ&���׭���:z[,��EX� -�8\+X3?�`+Kk֨���-s6?�dX<YIR����((�*]�s���Fo�IQ��(A�Pի�����mvl�K>PS� fG���(�\檐L�ƘԤB�-,F×���o��������Y�*=.	�c#�*%���X(���`,1�M�-�P$�VZlSTcM�#��G���X8*��L���R��D�A�i�_i�4�(���]!�2�نU��-����\�9�B�T�H[��ۊh��~�)���v������M�$��8����Լ�'�x��Ws�f9��!<
�Wv��e"DQ�47#ղb"2k�6�$X��JQZ[�[����y_���D�\�u���]��`<iE\}_+��bJ� >֏�0_P�Q�L���4=�e�$�#�WC�J���Ћ��>A��>j;�{8\����Ƚ����|�&���BI��ϓ��YOO7�����[���z����e(�,�&&�̗���ժ'��,4�y?C����S;����U���J�[:�+۶�Ha	U�m5��2���t���D�,s{JP]����I�0����i�94��K��	)�������掴--,H!��E��a��E�S�J����Xm�'w�%��Vlz(��ǒ�����&
�Zb)>W����#��/���IϵN+�;�j��K�$;��K���S\�\Il��ʝ��בc�R#������E����!a��Ƃ��t*%���z�
5�]�]�l�ᄏ�q�Qp\)�pEڤ���2�|�F���C#TW��O����f1Z���)A"j�r5�(�a��q���E�P~��A!��Z��F�VK+U
�|�_�ֈ��h���4��}?�g@Lj�c�9�}�B�f�s0��_o,Lw�o�N)x�S��׸P�	(�Q�A�V<����62���u~<�L������������lC�[VVOI�ȯ(ض��pRy+XfS\�`��
�h�|kW1���8��X5����4vLֈ�@qy��V�*�yp{ħ;x�ƚ4��(%Ift�?��'�^��S�`��y�% %�Ev���Ϝg4��9�fj�GV%H��O��(R��/�&��	�01�c��N��x���5�Fg�;$�@j,���ʆ�g}�]�6�:%ů(�?�3u���AA��A��--���^�Q0�&�YY~�γ�k�w"�]���^m�p7��a��$xx�<\�m��JA�B5�J�I�z���U<2r��`4P��,���?�75�h�����
Z���X[s�}�3�[\���Z��������׬��^����"�Uu����tL,��.M�A�ab�B,!�f�kO���8�� �33l����ljbF������v�����~�|֕H]���a%0k��~"�[������5�~GW' �h_J쑶��jV��	��ԈcX��Y/v�d]QG{��цnE��s%�3b���w�<�z}fy�4�,=KT����ki'p���/�ɘ�ř^�[��]	�T�%is3s��!�S�C �iC����T��Ԋ���ە��D�I�%'�=!��Ԗ�|v�&Ff\*��3!.�?�h+d���u���� E�bk%2�OX��۲��h��Z4+�`a��B�mxB#��!D��%��$d%6̉r׸�<�����L�BI�Z�RN����S{4NLs?�Qt@��7ht��$�ϖ�L\3�j�ZBJ�uh 
�1�yjD7\��I�rػ%~Mɧ�󷁝+V�ߍ�Uъ�5�3y����lFcx���W���PW����T�6K%�6p�]Q��^����k_�9�`�	�Ag��p����p��鄁k��8o��8ϊ�ߢ�k5�4�� �΃�ʓk��)����&�sA�P�3<�b�E���dLO��ui"�Sʄ쒨4Z�,X-°�'���FY�ZV�9��[��i���J�ܴ["�g��R:'-�#��(j a�������WF�2��B@1���'�:a���4�[�3匋�Ȫ!022:�L�r#6���D3�?�Ac�v�6p����Ғ3	�t1�s��N�G4��J6�?;���/�J=��T�^�M�/H�����S�JRZT.�-���:���=�t>��M--���)�UVN�S���_�{(;	�� `�|U*���*�q�H�MHJ��$�.�̑XX�b��xA<��A)v�pQ<$e)
Vۋ�c�Bn��LV#�1���b�๐�����h��E�a�3�3)� ZY����J�.��vW��@�Eۍu�rM�PƕQ�>�������`�uv&�ɯ��a�v��vY���|}QeՒ��?�wv���΅����`{��M��4�"�40dkwӒ��@ r�\��!�-&�}kԠ�LWG��bF"�N���0�o�;"�����u@�����+��/q�5J����Y[�?����!0�[�s/夥t�`X��� �;�i#Ҵ,��c-�ш��]1�͎�mH�� �����^��-����&�g�'X�M�b��ޔݿ��J���Lِ�-f�yUB5��}�g̾�ŗ|'ɂ��O��,��c�u  l~��,x*Ew��;u��l��r�e��L۰� ��E=SL(e��)���#1�0���˺�wsH ������Ĭ]~����|7 >�F�<��9�?c�s�E0D���%E�px&�Ax]p�=.	���,n�a!���F��u�uX������Hcz2�����7#�wh �>�B���Y�)*Y����n�t��h;��ӓ3<��^~�s{DH�:Sv�`���U�̓[]�<5�u�����z� -�!g1|IZ�mk�;�a(���Ru4,S�6����"D�h�$�J1l�(����l���q��?Җ�\"6L��hr%e���H��dQ`�w�ǜ��+�b>�ՙ<=FLO	�U����h� �o��_�&�i����I[_�t�,%k�D�ϻ�g�+I�%k�b��C %��C�U�9�Qh[��Q�P�?��r��աpN�(��N4������X8[!(�"%%�lm��8m����z�%,�+j�����n~xE��
2T��Q(m�ָ�w���/�w������
Y~���Cv�uB�%1V9pV�Cڊ�?	X �I�c���aK�G
�� �_m��"R�s���_�����X8�aU��\^�Y�,��d�\Y�G �&B�c�<A1B�2	�vp�V��:��3�V�R���I��I)Gtf�ݹ9&z��B�}�A�ř����-%�ҒR�pk���O�"Ad���H����'���-}0�A�d���_���9F��KJS�ق:]]�@�YiE�[�k�EuX?0�o�A��`:Y�(���6|M~� Z���Ҳ0�I�(;x�ؒ���.":�{H�2�L�Atr�KW&�'��KhÑ�[��>i�Y�֎eN��dBΗ :��{����A�W�EO��b9���ج�ZQVcI�J�\�(�
N�Z,�-�%�%����$=��q�~сI��4��_= ���^j�)�'aջ,���!\n3Cs>��ڏ���Tq9���¯��?�킽�q�G��U{���&�[B�e�"�=�*˿nٙ5���>)&��bK�����|^���̊��=���p�o���ҍ%�]�oPe�2&���%�y��9�W�勫^�o�>�B�������t/B�䰒�DĢ�8r�9��5�"�� e��Q2=e�6�"��Բ�_1VkM� �#	cMcM*W$������mmq����Yr���BdtȢ�Գ�H��7&�I�z}MB���M� �ҩ��W>������j���4�^$:�&k��Ѥ��;��8bBi3��H^�Bœj�13���!���|E4��/%�����Z�H�x��PA��4���6h%��ѤN!�ia�� ��e-y5��,����%I�N���}<� b  ��3Y�Zal��0��Ay��˧JJ��2�S��_�I����ɥ�-_=M�ފ����G��银�ZWB$&A���c�
B������D�I�⬰e=yZ���[���}�.-�ϔş+8��eP�i���KY�ڑ��?�}�SOʢV�C����o��I������ ��B��[��y�qc���-^% �∬0�!��"G�d�(�pZ���LV���D;t�u�n�>�'3��_N�͖���N���,�Ŀ�O �N�y��O�9X�k\Qz '�CR]���-��J}f?���9	�A��jT((���&����r?��HͣFJ*w_�5��.��d7ջУ���Úec���vɕ~z�g_yyo�����uY���]�jK�;�{�k���%��? �!��\ú:O@���
�c�֝�`W�%������e1`� ;�ǚ9���4���h�a�8q#�� �ǜ�]���Ȳ4)>��*��0찃�0������.��FvG8Z/����yg0��h�X\��4z1O�.�+�c^+����	Z�7+����K?�y��O~ʙ��m�ni |�5�����$O`��}�2Q�bvv���?�7�`hX0���ǖu=��J���'��W�7����y�t"��,#�`9�1�S�z`�! �̇���r�Z*_�ґ,�����B����c�;�2�A�`nN��Wf ��,�)����NUb@v9�0�څ_Ž����U0Fo%��g��8WP�j��9��o��0�d�_JJ���ɉ��B�=)	%���!1�����2��2"5R�{eAI�����(��2%��x���ZC���W^�|8��4X^�sg�(�(I��Nf=u0p^�����X�� �6�����ت|0p*�}�\�4H�]��Ϊ:��k� 
�������@ r����Y��{*-Ik�A!Նrˁ�a53%$�H�?�Sh�p��:{Z<@�F�07���\����TV�^�f�ip� (�Yʩ�yiaYj=����f�f�,A(���I0#br�S�?�c�c?��3+ڛ>��E����*T��d ��?�&�;3?o����5��K�O�,Y���j��I*�E. 0X�DBW-؎L�����#D��LB?�dE�֨/0��⒬k��P�U�섽0o^ȑ3���Z����@p��1��]�g�G`!ۑ�X���Č,��i�֚;����]Q�M��Y�/�u���g,7$��+�f�B
�䱤N��*�P
##"Y�����r'���4���X$���~��^/Q��c�[|��F�������cQ�NtbuA��B�=�-<WQ��e�B@������������9���`8�Np��=�|�$ rN���is��6?�����k�Hz*��Ȍ�A iH�N�VY��t�c�q.�$$bw1*�aX��na����8G#�֫��a��p~s{RVmC>Ǌ8x0����`�[7�E}ú�vIa(V��@*G����Y+�HDĔ`mK{�n_aK��Ͷj���O�W~�%4(�E���TU�qN<�nkw������C�RthH������������,D]���o�/�ˎ���u{���ʊ 	�*Y�����[TJ�����I��rc{���-ўw��������wd�rb�u!A��}������vC/�yt̿נ�>F������wX���l�j~�b�5ag�H2&�������S!��_l��r%G�؅L�r"����0c�qc��������������2��w��F+H)όgA�d0X����{�t����U��}S3�k�x__�����$`�L���1 �����}�~���>����=����za�O��I�a<��>c`	0�dS3���ESQ1H����������%J�h�x=?'�����ċ: 0�'k���P��XB�vT���S��N;��AI&|��}A>��H��
A�O@�)m����0B�.bp�u�Y��@�O$XqP&�LR2�f�</���R�li�;m��[_W�-�/���o����e��%d˯�mY��t����o���|VI`�G�b6�M��Ϸ[�%�?��߱���Z��*����K���OQ���¦����Ed��3ٶU�,~�
�0I�z�Ξ^�?�%�U����]z������Y"��1�.(!h�#�%C�x���6J��᣾C8��5�X3�7�����~�d�����p��Y%<�����G�эP�|�WV4��6��1ABi�(�!W"�(H.㱸���h�N�LZ�dU4X�`	��Br_²b-�l��$�k����
>�����|�J���脭���{���
�k0f;_#����H�,�����74<��2�&�F���1�<�%2��M�o�pM[g����° goyq�إ��Y�b-JP���me2����F6*��a���ZN4&�X/Ƌ��&݉%*EAQ��p�l�K,�����`�y]0��+9Ԭ�)�Z�!���Ɔ	Q" $L���N,���!p2繏(����Lg�Ji�YKW�%����<������=i�o�D�T��}����O��MM��̔�/
n�ӭ�0D��J���GR�`0I�.d=�Z��Xm�ߕ�bG��7����گ���C��g�iC�{U����!;y�t�߁?�<5���좥Rq�7J��u\�F�R�����׿�����=�B� A#~���q^�Y����]�-��dm$t�'!�R?Lnp��{Y^ұ8`���D@I|����ߙqpT$��|y�)4A�<Q���>GӍ�0���O�b�Fk�d�LIc$A[���$Z���׊iC��|���1�]`�:��V�⠌�E8��9L��U��e%�~�+p���W�$����C[�CB�z0�4$mY�../�>�:B�+7�{(��(�kɿ�r- "�8�H���[I�G���b����nrW���y�����F���h}XL�Ǖ-]U[f	�5b�0��#	���X�Y�z�ƍ�9S,@�]�TN�M_E� � $3�3������V�s��"ض�8/��'!���5V�Xcm�µ�R.(� I�l�;%�'X���j�%�|���[���Ξ>b#wG�ܹ#B���Oa����KP��	$�"i^V�@�:��@*�BƗ ��ؤ���R�^��_X���1h��}K�E3��s����g?7�BЈ���Mi@rXk�s��s���7���OpM��=pH+�|�=����R�Ї�L��z�)o�Ø|f���(i@��#9�d�/HPIN�27ʗMHQ-��S GN�YK3U����]xX�\/�*נ�6Zm��?0�j�ʾj?4����pb�q,ٵ��� ܼ�%�U��jkKXkkD�
6:J�4�:�HD�p"�lI5س�ϳ��΃z��֐��A���߬Kc�_m�y�d��%Ar-�/%���T�"��)ь��D��t�$��Y�X�@[6w$'X�Q���e����f�m�Q�c]�oC���Û���ۼgg�˭�y���+�3-�H�����IS��oN�[s���a���E/bt�|�xZʫݮ�Şz��0?� ą��e��ݽ�z.t���:˪ߕA�F���(q�����~�C�RD�3ܚhPs���ǟ�ű���R�r���h(d�zj�v xW�4jJlEBGy�FjcrK�&P��8���X��<�ZB���&�J�D~3%�!����%+���F��̧�k{��G$Z���K�R#���Z�EÞ�O @���1��#��D�j	uo<R=BS�I�`�bff�2s�y��z��aM h�޻�p![��R��^]�������QdP$���	L�7��|��V�:&}qa�f���4Q�K�O8����E�|� �G��y�!@(����;`|��h�WòI��P�A��c$�[�>`��F`�����:��|�d:����#�����{K[���{�A��p3azlV�p��dyұZ����v$�����:;���F�Sm-�2KɊ�+KV%+U!ǿR�B�"�Pc��]K�o[��dњU�T�Z�\�t��A��S}7��e�}v����g�p�͑YX��_�楤$���y�2h�b�z]����!��Dj�H�2��8\$��l��SЍ�!9��g��A�@X!�"}��!Z�C�Asa�y�	��`���eaY>D��I[�&�����cd�;�pɮ�k��o�����!�U�7��eV�4���<���<Z�7�ٶ,R�-6���b�����I�*�}�w�9��M�Kc�-��5'}���1�������u��g�Ia�Td�D����_]��!�bP�K�ܪ�f"3]�iK�
9iNY>j�1ǀ�eM� Y�aK�5�>�D@-P&��Tc�ؖ:��qU�B" �WXjA�J���^+�������j	B�5cNP��%�n��/V�"������C��se��#Յ~�5���z)�a�����G�.47�mY��:52k%�{��[{b�~�S]�^�������$$�������./X�r�j+�R�)t�3��JK�v�9�g�Ȏ5��$���뜪=��Y�Lv��˭���:�����7����� 3�_X_�щq��v��!��sg������K��Mcf�<<?3m�ܷ%)5,H`w�e.�˗��z8������(Rأ�+��V���(G�;֐\�&	�ɽLA0H,��VJ7C���Q]I���9��w��7���y��]�F�L��9�-��ø�ޑd	Ҽ"�z�����N9>�?�q��z�lN9�eqiWg�Z�664mCw'm�r��X�\���^e=X�.0n�?���=�1&y77W}�T�I�U�pBˑ��A*0��7
� D�� b��'��mA������<;�!��v+D�������&h�V�Yó�Ytk��>Y�̛Qc��c� ����1��2݇�f�64lfv��8�D��f2b�--g��U�#d]]8��6'�[SY��'�/"Q���
���Xf��J0�t����ϟ�֦:�@yT�\R4��Lh���H#����G>���h�z̝_X��/�mj#n����>cOȂ������W���(X�r��T�u�������GCv���j@��G�F<R�%�&�v��y��n1����ۥK�����vg���5�h��G��B	r_���PԻ���a~���Mã>�?����3���b��#I�!���_�7�v�X] >��7�l��ƃ��1ڒ�nZk[JWe��5)e�OĚCrc�%?�ĸnZ�PJ(��F���]��"af2��c�*����%��m���*'���:�c�(�`�G�P�!���B����W�'?���s!-6VY��{&��@(" �J0Fq�����%�LJ��!�=��n�G���7��D�����+a��z! �73��Y5��Z���.u�������,��jT���B0&>A0tNV��v1Q�����'3�$3�A g<*X�t�s��ta�%Y�c����@A�@(�Z�֎v��o��c�� G����G�o�5=O���"�2`P	!�'�8����0}�KE��J�FM�5��ۑ���o�?���<�g�lnf���]Y��oO�^�R��A s�Ѿң^�sF#q���ՊP�ba�6�XIL��%���[H'���|P���0w�O��YJ�#}�o��7��;�>�9��-_���`�B�F�,��K�j�V��`Ѭ�u�Y��>�������:r���|b�q���ŷB��X��	����%��UA� `�(oe�gy����B 7,yH4���Zb�q�k�K�H6wC�����m�ߎ���K\�5(z�WU8t���L�Mc��� �tb5pR>XX7 �����t� �F�L<%�E�2��#�D���`�芬���1�����-$�B�:i�}XF��L�#D�.@D�0�ߤZ�F��6U'`�03�d��Y��`,��Gt��*�d7��j�s�FH����ʳD��;r�={�|��":���.l���� zoy�I�"��R�1����ĞÈRH:�y���lڭ{R.��5�W|�?����}��e�}�MN���ؤML��Җm�n؆,s��,Ez��V�Z�b�&c�����[ِ[5�D 6�gd� �F��1�W�A��_�g��(b}��\�BU�=4&��*T@�7�(�����nm3��Ҳ$1�bQ�V(3�0*�Y��a≘%�lYN��%]js/�$�Muߒ�"�#��FBv��D@o��	���s%!�a
��Mc_6��t)ؙjik�A6�����g�#�ˑ�"�ȫ���,��-m'�MP-�B1>(��<�7q �n���E�?�ըc�(����8~ZN3���3�X R~`1��SZ�pY�|.dR1,�5�&d��Y�)�p�?e�eI�=C1�2K�$�� �N���,o����CC6��}�Or���MM���6M�'Z	hK�7Ұg�J��t+XO�4;�<�9k�j��?@x�̂TΠ�t��h}�7�ͳ�&�mlV�����:z��@����KҐY�iMBS�κ�|�h�O��I� uQh5"��@���UV'�i���[��P&���)�-��Ax_�C h���3��`&�[���4��ch�F9��s	�Y�ܪɪ�b�����g����=l-�R�M^^%��&^R�@>d�P㰭�َ�p&mhp�!�,:YzE4�`
V��H�B���h�h"�A
�2$Hlk��wA��s ����-�4x��$���9�.Xz�D��l���F�k�V��=���;�:��b�蕘��xl�
I�s��j B�s"(,�j~H��a���7#�_��Z2���w:u0��/���h���5ș�ƪ��`C� )AB+���g `�� dZ&�&����)Y�%�Qq�����/�I�+���Y�M��΁� �,`L��{�Ũ�>�b�)�sW���u� �/P�(YU׊в ��^���8��!��Ps��߱��e[\޴b���=����{� ���+����֗ڈ�����"K�ei��+���JNV#�/�m�0��n)3]��]�,4-��jj�&�����5��+��R�G�@�<�E�*�{1��)_
�Vc���jO�I�����OK�<qĺ:��!Xk*�6;;�{�Yg{�ܑN�X4a[�奜W��w���feɃ6�?�)��(~"��յ�[��Gery֘�@{��L�2Y2���}E��9x�њxV��=-�TXD<z�p����X\�9��;o�q���}�)��*��<h@aO�."J0�Ð=�|�#K�7�!g�!_)��{�G��`��%Z���aS��`���	Q�K"�00ͬ��4�4u刟��^�`M�ͫ���YڅB�����z&"�8 �L8���`
u�����(u#%��l7�_}��6ss�,���H�a@�4D��*iHiXy'�_`�x�dV_�U�e��k��+�f�^#���LH`��)h@idk�Vؑ�i��?\__q�0��=����]pv�I�%B��+)�v��b ��gR΍3L� A;�*�s������d��ȟ#s�����hLg���{��|��G}tk���q�O��ؑ���9;4�m�x�#��� ����OCɽx,!��bO?���E�ċ/������~[������#_��3�R�G��ecc�p�m]�U�[c���Q�
4p�.����@��Av��j�U���Y_S[/�J��W��S���ݨ�rq�d	��|0���"2|Ix�0/��h�1EeE�N�>m?��س�Xoo��^\S��ab4�B��,Y�켣'�!���QJ@�"ABX+}naM�5��j�i���1!bw��
GryqŧH�b�?B�,(X#��LBoI�wU6E�|n��u"@m����m_m��(�H��M�a��rY���ՆE��&A�z10�F�Z�A�u��[����
�N�W�.ЎP�/���I!��I� �߲��Zr�L�bѨ�>5)k�M|���&��CƼ�[�c�Ma�!HYh�����Р��׬�.�֮��j��g���t
��%�Gl(H����c����D�2)OYm��0<5�۰�^W���?B�?���7Zכ�3l�L�[�0��?�����3���b�Ը�9J` �N�&�<9�{j�0}@��<x�	S����	� �C>�����;M�3є�j���������X��A,Y�t�Q7F�]1�~�}��A)<d�� ڏbb��Lh�E�R��'Ɗ��mBc�H��X_o��9u��[�퓟|ھ��g��+�KW�*P�]��86�僸^�R�����	�K�����pMO���R��2�?BɤrU�٥�=b��am�)~���;Ru!K6���u��^���� �aq�I�(� �Geq�j�:7d�5,o��!K4�ؑ����s���9i׳����v��y;���v��'��c�}�'��έM����o�+(�)v՛��,�3�UK�#OQ�^�GXV���"���BzHXo��TV�a�"�_QgB��
���k��3�*ݜ�f��m1
�1a=�[�����1�P���:����o`V������az���>��kg��,�~^jlξ��{w�SQ �E��ח,����N�!4!�b�'��z��MaZ�#@A�}�EY!H(~�
*�,��7&r�cL�C0�Q�,���X��弄e������7�
����߻i���=��r����a�ϡ�Х�>���� 	����R�?)�4ot�J�l���7�|���(˅��������XE�`�ədv�
	�� �B3dr o�;dޭΓ}�aҞ��dR������,l�(wH�T	VI�cIkH�,.M&,�H�Ye��.1z�7h�?Ъk��-���f/��}�_�'�8.Xr֞z�=��I{��9{�ٳ���g�iA�ǟ9eg/���Н;v�H�z�Ȼ�h�|��E� ���B�|�z���``�5�w����p݅�R�����	�Fm�R��ޛʗ��L����\�L��(��,����p��@P�`��P�^�	Ǳ��#Z�/]��La� �<�G���`48Ȇ��)���ͽ8�2)�ɔ>~����e�@	��,Ya�Z�l�L�)�@^a]�Q��ʬM�NXU�e�K�YXqa!��c]�}�j� ߖ)��C �����x��(F�μ�D�	r���$0��L۵�wl�ި �|�U��Q��H	�(��(f˸H��:7�lTE���e*E(ڈ�nr��-�	ζݸrݾ���V�5��8�8�hL$��`�:	m,!(VOCIH|�0y��.�[��|
lRӁĕ%v�tR�ٲ�3���WU�`��N����ӟ�3����O���s�# �퉧���);��i{����s���~Z��3����?������*���s�ü#v),�|E,ڊ�+q����t���^�G�����a(��$�|>��&�w�n $�uYX�6NTlvjA����Pyx~~]�@�֫�Z�콷/Y.S�� E8�V�O�ճ��[ ��WI!�%���~�G�H�ƏBVYbO��gtƂ��-O���(ܔ�����گ*;�J ���"��7s�G���@��F�!���D��qG*%dmR�Qo��ϙ�i������h�b]��_�4%�LDQ�%��ܠ ���1�J(��&�l�#d�T,��~��7>)��`]>j����ԯ�F�F
��れ�Q���E�Gj���C�f��,��.
�9TC #��8V�2������_{ӆF2�R����H-�k�8�0 ��P�	�`{�f���b�8��6-�/#�
���N�L,���K#(�m��5�)���?}�������ܲ�K�_�@��2�,������ -�x��T<nmM1_W�_���;7��Տ�ڍ�,#"2�s��]�u�]�vϋ��d��kMm�уT�
������ȷ,���;Y/hպ�
c�����p�a�8�+��s����hQKw؝��4.�X�H8�1l7��]�����kC�M��u,��w�|��:��5HF���T�����X i��P�y��9��{� ��W�XG���
ƞ�$N��!�D2f}�����O��y�y�>��K���2��3�Vf]��ԣ��$e�'�&E�2���-�s^$�[�>*�$�c-���W�u�Wro�|,9�L���~�#,�n�L��4�qъ	r�7��C�	���-ʭ��~��W�ap'ɒD� )�ߓ�%9�`�>x����-{A2���>,���I=F���/��6<���"cDl�XՌ�a�,�
Y݋5*�d*!"7GG%�2��TJ�(�[���q���_���J8��L��?�j]�a��Ԓ�w,L��_׆F���]����Ͷ�>w�n߻#A�d]}�v��CN\1����9�t�:��/��{������p_�B=���%@hHˬ��b:������,�v9��t���_��y_�JUqk�����^̧��Iо�b�\)Y���6K5'��nM
���>�Ln`KSʚ�Ikmm��NYA���6��� 
�	a���~x��ɭ�>�hy�^�A�b�
f� &S���^D���-:t����F��V
 �Iم�ҢC�R� ����*���E�(�J�-��'��v�<D�m�e%����I	�|L����#r	A�#�H�^C���Az��#��!1�d�{e�D �'(�s�PB�|�Q)t|<���Ry�L�x� U��C����'#�"S]"O�P�:��p2�c"LL���ifѿ�M��)ݼ�H�����/�=G��5�����D3N>sFh)` s^h~L4>�dM61��"��h�yv��a�~�q=IN���Z{����g~����g��/^��?g�uY[sĎϞ��?q�^��y��`�������Cv���w-��Ѥ�2rї- ��8�đS-���?��ض�8H��@����峾��"Q=�B>�6Xg����OX����-�$��LW����F~R��R��612��\|�1{�����=a/�����'/������G؁�1p�]б'� *?n�^|�.���{ʞ|���t��Ԭ�uvh��lz�}�-R��g)R \�L����=Z��5y�)fq.�:�(��|�/�uJ$�v�p�>t�Ĭ�Px��K������w�|�Y�0wu/�?#�C�7}h&SгAj�C��p���g�BW��T{�>Q�%-L���amH ��FA�/%&�`���ƤGDER�%$��,ݗ����H�ڱ�x��kyNy�@�V�������Kb�U�"�՜N�J8u�u	͆���ȇ�h�t�QG(��8�Y	���{�%9���.ՠ�A�g�y0���h�-������V�Y��i�*[���F�CdH�Æ$�-騵��$�,d��E[�dmQ���N�m��Oah����tnG[BB�c'���ѣ�V_�g����)�i��g�E���,�׼\��0����&���j �jH�`�� �L���g�gIL�0����b���?k_����	�2�bT���*1з'���G��o~ho}犽��-��_�c���7t�=���iU[�Bbr�$���R� mLO���dא��� 4A�rǵ9Jnv�S<�E���ч`�$�!P#>A�AM�ǘ�"	���x:�e�`���g�/H�g� )ݠ�(�εtpo�����k�s�;�2yH����*����r�śu�����ۖ��e��v��%�E�rAR3��yI`/�2�E��� O�yւ�4�d�T0�A���P�I%u�:�R�����D� Z*��0g��J��z=���h��F���D��`a��ki�r9�	�}�N|)����������}�*+���&k��v�S36>:a#�ldx�n�|`ׯ���Q�`�ɺp�G�쥗��W^��}�s/���v�@���d�#����L1���*�`�op��T[���Q����\oҿ��$N�(]ý��W-�&!|(yA�x��S1:��w�u_]��;�pF�EsG����:�{����Ko�~��ؔ9c�"�N ]� ��=n����c�����6��kܗ�� ��_~��uT�<� ��qh�B�a��c�ן~<]��;���배4��A)�
�D�!��~��>m�o�������N	���k�?�v ���;���`�։G5F\�3)zD�e���e��24%7���,#Bu,�{	�-��*c������j`��0I�>�F�^�bYқ[�B��uS�kf��֘�TR�b"��G���7-!��7�p��`4֍A ����wC�A�%k,�������<���$d�����Ţ��ږW������֖����H�ٕ�v��]�w�ݿ=(M�>|�C{���������G&|��eiwa����d��lh�ݿ{O�;bc��^u
��w��_��wl���O�����m��P�C`a(�#��*�cC1N=l���y�s���Ȃ�~�om�ɸ��k�X ����²}ϳ�����×>a������#�==-v����=�x�]:5�Nk�Μ9jǎ4v�a�ə�~<j������H��\��1g~��(bᘆ�Q�J0�&�ꅏy\x���`�1�f�y
�k�xf �%4:�}-�
|��@HȣZ���6�׆k��>��\�j�c���ݍo	��#0�H"��;rqt-���𫍏,>�SU+4 �(�8�r���n�ch%E���(G0rd����`��lfI�	�e�l��#$�@v��tXA��QZ4,YF�^<�x�\5j|���ypxIle���b9= Y�:��ܢ��R���{֟�n���KW}Y>k���Gu�3y�������,dm�jQ��EY���w���؂��ၕlv����ʕ��׿�����o~O�����$X+�RYi2Y	~�zQ>x?z9+��@jB��$a���1����򥬲�u�n0��c�Ǚ�ے�,�����PP��]�9�sK�7%8������ FV:��)�䀢��D|����R����&��B<g���8�yf>����f dX.�ƾ���~�a��&�c�j�k:�L��B�����_Ĕ���X#�� $���(9GFL�@�F��B��:��<�`�ݽ���ϣ�"*~ceծOd�EѬ��i�,�.�9�A�5|O6Ft�'���_�8&᜝]��E!�k'�����������K2�Y�ȼ&:��]��q[��I#	n��2)/���nѨ��@zN�P��(ɪ����g�,;Q0�@�u9l�N�F@U~ɲ���ߴ�q��f����v���i�����g.�'>�����ɏ���>~�>�����~�R�	�,e�ڵ����ٕ.K���\]���[�Z�	��j����k�&�V$u�t�.Oݏ���D.��WV=�U�d�<�$Bq1�hRY��fkE2*D{]��x�W¦��ZDx��	$ؘ��Rffw��.0���	l-����7Y0U �����,.�3�p�CRz��VP��7���m����۫1s+���f��?����B�7P������<�v"$D9�:JȠ?~��Y�.>.�QS�I�\�t̟��ҽ9�4���w��q���`��D�]�ғ�.CB�!{���dŘ�e����Ӷ0=�u�|��҂�!	\`��o��Gb��т)���_q*�ǂ?$�ac�k�:2x5��Wiy5Bme���r�e���gl��|���8R�{��hhƚ�i,{��FC#�@G�Cՠ%G�8�� ���[�l����`쪗���k���nu��eG�١�;6�k'����=6p�����������?�{�;�83�@hA��p�-��Vs�D���g�gx�|	Vy�Cڍ��d���ۺ�P�����id9d� DR�1��M��\=5M�( 4$��t�l�z�͌���ga&=�7��i�:/�G��q#q����� �#���"e��D�N�2��`�m�f5HJ&"]�ir��Q���	��o���i�ET�fRk�y�9x���I3#QkL#c�b=���x������wzs7,��7��Ad��7V��Smb��u�)��#���Yd�-5ge�r�ߔ��0�+�X*`��*Rj��d �XL��5"RF�;h08x#Vr6*_ffrV�Hk��������Y���>_���T���Z2 8�`{�\XJ�'���$|�ݴ�+cG_���V0�@����e�����^2P�Щ4�/F���3<�V�@S�	g 2���6�Єh��a$^��g�)�f�,�1�⛱.��b�]���l�sJ6���a���Ac�~h�������X\)zʙ��B`9cB�*S<�q&����7H |�쑰�O���9���c1�'����m�J�/��X�+@ #s�,�$��a���dp&���"�HM�֢�Cs�@��|�Lox!� ��s�� �ݪ�8V1�K&���~�x�f��:��i��c�Vܘ`�->f0����i�R�Za�	������,���5{poN�_r�k��6b�BpL@��Oǆo��i���=��2����-�Q��&@ i$�	m�����LL�+'+��>��H<��1�Mg�]i`��A�]�8�@V���-���}<�D�9aŀ\�Ҏ�`TA���a�і�	��!��^ʢ�rσ0`x:���j�O�S'��������K�I;p�ߎ?v�`R�A�fل|��m�����r;�H�з��vY��z����z9���YB�6��g3�65�e�r[ߩ���ˁe����H�X��b�:�R*��o���_�����k�W��z���Kv�꠽������?�������6<2i}p���/�k����6!��B�}-s��r!DR�
�1�1@ ..bT�Y`�u�<��~k����
�\=؟���+��F�F<�,��n�ynM�s�<~�k�E�_%����(�D��-˗x���P��a扬�����I��>Lu%�1��u��
9u��F6�L��	����M~�_���ՙ�%�>�����oIi��
/�^Q�Zd_�QxœFEp5|Χ�f�{i<�#�A��%�dy{�{9�8������׃��8'?�_��Vkv>�ZA��R}xy~�V��QM+;;o#�G�ޝ�7�&?�E�E���?�Ν?f������di��a&<Kv�sv��v��J���z���lu�t Y��W�(B��>olUӛ�
��ە|��<���v�����-+����/���R&l�$a;��I���		�q�X4��,��l��_�i��67?gCc�vo��g3TA>Aj_5])�%�����]�w~�=���VVV����f�D�&��Q���<���� ���:^�4�(/�N:�J4�d���~;x�W�a�<P���jv"�.B8mR|�+���g�����D[�9�N���X2,)n�,�e<�b���i(j/r�Z��j,��j��>y�
ód�w�%�W5�<	�<Q�Lń5a�}�t��~	���$_~��ŏ�Ð�/G�xMm��;"/,x���A�]b�O�EKbJo��LR���u��&�ub�1���AAsQ�Z�@�}��"��?׀��rsh�Y����܊Y��������6|�ݽg��lL�4���|���<,s>lc�Y�;��9;��QۖP0w�$��"��, ������u:����W_����	��x��Ѷe�$u�V;*iZ�?��M>�|��XD�'X�{�@�$0 �� �/�l�5�?��[}ܢM����]��޺j�~�]{�����x�C�y�]�F
ٴ�W
>�[^�)�#;��rA-�a��ڍ+7<M�(���e	Ura>q��eV
?�!�h��.`QB����%�9����	����#8F���xj���>��>\^��5h�@q�]S��]4�{s�d�j�CG�lz"cSS�g��'�?+��V����U߄0tP� �#1,V�F.#m��[�{ �o��M�})A�b'������*�n�dP��\&�>|:\q���W��r��zcKL`,"&�թ���ب��s�`5ֳb��v�貨o�Z;SM5�0�dW������
K�Ɉ�y����kT'q��VO� �p
���b�I�IG�,� H��l[ky��P{7��no؞:���;��"&���:lO��<��iK��s��8���M{��kv��gw�4:z{��#a���77w��@�:�BV�?�p��ڕUZg.O��kP��^�0�#��f����B��;C��y�si�oy}��S�������Gwlzz�<���q�$���²�\i)+�b�%R�\��l~.k�cS6+&]��X]+�<����@O���`�x�0X|]9���{Ў#
|��\��s-�U����a�DF���&q��a;xKFZHHVV�B�0;r��
.�֭m-�ԟ �����phHJ���٧`yUt��J&AC��my�ٙY�d��A-�?�<�J]}��.
�ﰬ�C|o�����wk[Z�\ƤV�_!�$��\~)prߪ��*�נe+�X���Ɗ�
K��-���.ʂE��`�u��-"�?\C�7au��߬�fcjt�!B���Z-�R�5�yCSi(�CAZG�]�3���.�Y�g� ��H����4-�Wq� &b��k+�AG�6�G�8�;E4�/$�n���:	9�mh'��Zmlj
[߁6�R���aA���6;t���뱄�	��`¾ �̔�g�˚JiK�V�5�gHq �����w�K�z{�jY>QS>X��)H>}�� �`�՛V2�4�;~�|ߥ)[,�ۊ�rOMF��ƚ`gQ0q���N/��mH�c��t�9C��y2�`8�ѨڌK�4�x?�Rj?/٧Tt5��B)��͸xVZ]��1qN�~�#c�_�?��ߩo��9����,|�BO=���ډ�Ab0�O�w�L���` ��w�M<Ƙ#TL�P��8�> ����^X�f�Q�1"���~�EeEc�F��te�Wg�mjO��ʝaE�X��:Z���%���X�A7�a"�Ma�&��'�]��4���Bjp����@`�a'�D��(F�{�G��K������� �.1��j]���]ח�z��<��a��д�IK������h-v�L��� �������uwE,¼PE�pA���E�
�mM��,?A=F/�\���2A��sd��]�	S�A���E6�RN��r���喊��cS�Y�=����L���ۓvx�{�����P�34����9�F�5�A��Oi�������mz�\�w���	�/���C �(<�������1C`8]������p�
N��o�8��֏��x��4���q��u/�O_<�C|��qմ��c��?�'�;q^����zq�[m�A4�C&EL}u�h�b1'Qg�wD���>��}�OyM�,7�R^D(㉨�J��`�Z�oah��V�)˾^����3�X,M�/I@l-Fh��W��Uvn%��_F��A�n���u
��3�#���t����Rj�ݪ\3�1'+�c@��E��}����|��Q�.h�W{x{�ͬ���C��ݛ����5g��޾f�[����e��2a�=�v��"]auϖs,�۱�գ�K�l6�Y���U��ݐ������=>������Z��#z�lhb����Éu�ʖ��ئ]��f��)J�	��3����)%d�>�4�[|��$pC���dI�feE�	ڂ`���#4�v~��zK+S6u�B�*=˃]z#Ll��!%�-�J�|/���9<�[?��h=W��?��F�Fi���,�d��^��5n<��i���~���??���7ڍ�Fh�;x�v×�A`%��iA�Zэd
���I �p�ޘ�=yr����>mm���T�9ݟ� ����^R�2��!�-�,I��grI̳�YmG��g����nܥNa5�ո`y�t�J��ND��3�>�z�[�@�I��;8|�7ڇ?�:>_�`/�9�e2>���c� q���ߺ�K�%�@�-���*K�)���W.��?�	��Oʞ��s�jﷶ�C��=��'��?���:7���<c}��rU6�\ocs�:Uvwl��l�Ќ��l�ݟܵ3�6�Ta��+�ŬT���mV�lj�Z�V��t��T��B�͛=�-��)�=�S�`����s�kA�
�}R������>��F!��I1 H>�#���?�w�����7�u�G���\�A��;w�B���qa�R�LU{h���#x&c
���g�
�O`��j�7H��
���̀�<�,Fq(H[� 2"P��y.��ǟ�����N���u���	�1�<�B���8��(��`U�@��_�'�y�K���g5zt���ʺTy>�vBּ��"[�l��);��I��l`_��E;$_F&��)����~s`�}���"�\�$τ"���ш�P`p�O.���k8�p�*�l�F����.q��	F���F�7f�ٖ��U��gFD��)�Ą2;�n��KCb�yi�Z�Gbv�o�:ںdmV儛��y�'���Ŗ&�v�W]�n�Vؚ%�����F�,�g�m	�j�ͭGl��h#�*�*��}�q�%;|��,~�U�Ymj�
�1[/O�f�ޕI[+� VŬ.�b�nkP�����׿g3�sƎ'�,�D�@AJ�CCiz6���t��\��~^�ԗ���:/x��l��K��^�CVW��i����b����K��p�>~/���M�l} *���o����>���] ��^�1��h�3��o�L�?>ڿ?�F�S��ЏS�>�;:-�1 r<Ad��z����JVV�<?�����(���z��j��Ç^]�/�ґ�yR�,��~��7k�#����E,6,����A������S�w�@�z�k�O�LG�@h)p=��A,�V��c\�6cp�'��I1N*�(�~@��!2�i5�ư��C��MV[}<�w�j�6�bJ%��	gϹS�DpV׏�ڻo}`���}�[?�7^�^��7�[�}{��o������������o~Ǯ^�!��v5�_���Aq՚:�-��kk��ܕ�c�V]�R�]v��9k��sA߭
	r��r)��4ojo�������G��!ö��{J%טT��E�z6��a�Pp0!�_��vb}8���0����6�;���fa��� �0�7���HC��z��Ue=@
�	bDh�p��	t �<?x���5J���,.ZONX~q�w�A�[Z��httk]�\�MON[G{�M��x��)DGavx�B���h���@1�S�i��$��5/�
僕_έ8P"D�x�q+�*��w�wf�q�=|8a��9�'Qph�&)��:ǲ�_yyo���;կ�DE���K`d������Ea�<g��{n�ټ�b���_�UV���d��N"�#��BQ�tk��m%�H��#1���N�����Aߑ�ʄ,�v  ��IDATr��� �t���R�Ƨ"LM�y�:���a������gN�<|3�hDډDOB�붼8o�?�n���zƖM�-�fiK����u�,�k��3��4�L(�G�I0�Άkn��;������-W`��-Ք�-��1o/��@�Pؕe~>��,��@LT̗J�,"gyfl����}�u�ÖMix_�.�F�yN� @��M�a B�\��`4P�^��Q�XQ@�6��+V�+�Jy_���ߕ�ڈ��Z)�ĘY��t>_.�I��S��+M?��ܗI݌�b8p��.<���oVG#�,���l>k�$��� �755I�6���(�g�5�+��n���f���MQ&�:�~�_�a������@� �&I��Ew�ˤ�A7TKV�E+�]Pcq��Ɉ�������+���s��
��+�	�Ԟ,Y�����f3+�$;�d
�bN&mjS���-؍+�lnf�'=��}�,�.����aI��ym{��4B�"S;�syzec�����9h�@HР$.��m�0�hҚ��G,�NYKk��8y̎+��1�ԿC[����ձ�G3gg��ʥ�b"1@��H�uOf���[A	��zV��8��|��c7�t�F$M��ʢʒ�v*t%b1{��D˰����z��Z��i2�0��~&�	ߤ0[2���O2���V���w�آ�;����M�ш���g+�mP[�
,��w�V���|����c[�D���X�n\Jց�BA�+,##(��d�>&�k�����_-Xp����~�o���S �>c��$%L���)���ص���굛v�����4˛r"�SSs61�s��s��~MNֆ�lw�<��b�]���;m���S���;�.�~$p���`>�d�@!3�(#,ʃM#�=�^�ě[�OHQi�S�m��4 0�]Q�%+���_�.�H�Q7i�$B��ḟG�mfa�f��B4���z0ꍥX?��h��I1�H}u���ڌ(��V���E�po8�n��r:!E;U�ɩ[���z���Sje�e�Sc}���ӕv[�s�a�q�q�! ֍����w'l]���x�[d&t!<�|0�`�f`a�<j=}�63*�_���ښ����'G�Zp��g���D|qdTB�֌ȧ�����j��!	BB�w��C�XV+J jrb�~�����.
�n�@$SI�����6A���G�Ҳ�--i�K����f�bF"Zڑ���b���á������gs�=Q���>��@�	ƄI>��(7A���� ȅ���:+���q�E�{H)l c����s��[��D+BK,^)���>iaj��ސ5�$/x���̂�IH�r��@=wu4vX_�Cd� �?���45Q�/���Ge��<��E��Akg�#��ҪCu�i��Y%e��cj�ʁ�0l8�h���W�� M���z�YD|��~��Fl"��r����ma}��XAOc?<G�JH�Tgb��{Q���a����4��'��J��Mt���O�ŏ_���i�K�6��b��$�,�� �dP�İ�4�b챑q���Mi��_����]������o��V�
�����/ڳϜ���i	٦u��ؗ��=��y����m�0����8cS�6rҦ�2��ބ=��q	(��}������K�i{����[�wF�ݔ]V{�^�!%���"��"�=��ȑ#v��)�^Y��ϫ�W}����k�b�Fu��V[b|��ŭ���Y�������I����Z�� L�p6
���u�H�t�R���q~p�8 zK�yU��^���;̍ߒ/|:��e4K+<	�,���	��f�jt4��Uc��/��C�h7���|lk���9�?����YF ��)��P��p��y�<?�~��ȁg��[HqP�`�WҳA*�Y��O��wpV���C%���*�f�wuC19ЈF���H�����"��3�"�Z!�#(TCh)���cN�Ch� !	4�sq�,v�3�"��D��n��Sv��9{�c���3�����$��L��[�|���%�P��Ku���h/�SW���u�PY��c����g���A�����V�r��@VU�}�.~����/�dG��|�������dlK4x���%�W����C������v�|b����W��d�iU�(f8��D��,f�Q2f�+K.�q����W���^z�!"��^�}�m�	zr�����I�)�iH�,��5��d9�>��S3��[o����#u�Y 5AP�A�A�P�ҥb.`);����B_)�p��'~!�R~\q]�g��H�Ju��@9��!(��@H���z�����(L�ڎ�ݷ��uߊA�P���{�F����wme�ղ�PMz+&��+��.��%w����7��7(>$e����݈���=0����s�!d>�l��A��O��ɽ�� ���H+H!�'��0�:��#8�R%:����i����D#�"�X�uS$�r�%_�CB1��X*ą�Ae��R0F�*�ƚa)����a?���OY�U��"4vsaf���O_�
YB��+8� a�(x"͸��q��r�7Wly~�Z�������؝W�����a����U�T�t���/���O}�"7�1��fs���8�%�3o�Һ��y9�_��/H	�?*!��3�0�:�H���j�W��,�幄ߥ#D�ZA�y{��?�o��w��w����~�_�O}�9�y�袠eA����;v��a�\hh,VGVLHclbN���!i����D4&K�y��koط���MML�c�p�?���g��l�G�<j#qC �U�Rn���!�{���酐Ms�ZY�*����!��?��r��@�84Bi��4_�M�:��bEc�}C��g=��Q�;.Ae����a/=ր��i������HŞϏQŏ��v�](�;���K!��w�v��Rx�`E�,ȗ�{��l
�_\q��W��M7��ّ�M�B�A���@8�?�7��M�S��A�#�V��X��քp�;���Ķ�
���jBD����h@�I�ḅ��P�&���5��mκ�1�0*8T-f
Ym(� d�~ ��گ�C=���b�Gz���ݶ�Ҙ{5����-�����!��%�u�e��jfo ��+l9��Q�^�{����^���fkI�}�lO�{OW���v˷���@^�-�kh0�x)D,�*��j	���Z�J�.��jd�e}:�;��~�Ǥd"��8��aԬ4o�kL�� ��;�V:��U�A�T��,�]��Ș Zޙ��ﭱ\��/�3cG�קx���@�tG���/h��@���3��_�҃Ĩ@��� N�q��������c�ؘ�k���E^R�z6�ni��b--b�ku��'��p��Z	��X"�_^�J/|8`.�𜈔;Y�@Bwud���$�F���Q��� ���?Xr�a��_����|
=������ev����c �2�Wې�����5�*f��v� ��G��P�P��&�[�(@Ӯl�����H����c��Y���,���Oڧ���}��'����_ڡ�'쥏��?��?�;wرv�d��L�ި�>���!vm� �"Tm!i�w�}�-گ��߱+�~h���}U������ �����>���%�_�ÿ�Z��gN[�mh��Y>�����&f�`@l��nl�N��wD��|ÄҨ�����a�����Fʬ���o��%�	LI}��=�-9�y㡝=wD�Hin�a;�P��S�n��D9m��
*`��,�낚���=�Q�K斎'`ͤ����QB]G��2@[�s6���B ���<#C_�L(P��9%
��$�/�h�����C��� �qa�^��H@4��Iz.� /`�Rgw�/Hׅ%�A��>x@�)v֙a����u�R���X�U�!�Ρ��v������x�b��r��]^>�h0&����˕�V>�*��LcF[Z�A}z���.wI+۾��9�Ϟ�@`I���/�R9U��Ѥf\�γ��t�8��R�� �:��ށ��yS���l��,�X��Ā�B�� �����a�k�+��������'�V��ؔP	&�;c,�A����h]� ���2K���$���xCN��;�K��|��8���,��������e��BA�/.y���޿l���������>62j�c��?&�WM��&��1،� ��������L�����)����Yթ�q}����E�k��.ƫ����O̂��\��J��]�@O�i-�%x@IO��XՐ#a@4��461c��O����*�s
��r�u�1tf��G �7J8h�_���1,J�.��a��*��r	M�{�p.A�!�ZLa��޴uu��9���'�N3�M��-Bk{�WX�&�>
,ذ��Ș~@�PH<� 	>m$�?7��s��X$&�5(3�*i6� ���:��%'d:a�x!���}���ll�W^�&}�67� (%��3Ј8|X�J=���!�O����-��}P�B��+���g���: �/]�I��X:���v��0��f)Au�Uw�6%`�b�X���pʎ�%1}~}�J�@Y���EO�eӽ��u�I���umH�a�qSVgd�bMM�����Q{���="�����2h�-Y��,FAP�%^̑�b�C(�O?�d�3�:�k����tl�}�ʶ��4�Ѐ� &���1YS6⣿0�N�WI�D�3/?/����yy.5�Y�j`B%�N���#�����і�?X	��ʅ��ݽ{OPy�S�"0�����J�I[x���Å!@��N	�� :zo��_���V�EI�o$`�5w!�fbz�px.L�ps��=�v`�M���c��X!���iM�O�3��Q��	d�y��y�T�</֛H�$t5Xg*U�8s�ڻ�v�`��#I�SzC4�������$�o�X���fq2q�4�g�g����ѡ��\�o���}1au����L�椬ٺo[�T,�e�	Y���T U��i��SR�@�kh�#2F��cW�Qn �IF�v�)!�����,��M��f��wjjB���`_��?n�o~�3�s�C�!8�&�|�/B�:o��Otzz�|�Q���w�����￱m17�
D����k,�q���*�	u� �� �Ƥ6~��{�f2���3����=}���$>�=0,��@�S������N�������a���\*�؟�ٷ,��,l�2�D�k�Y�Zes��}*���t�hQoMɴ�W��ɂ߸u�&���ī���Q��5F,ޅ���~@��13P�m,X����>�ӯ!+?;�q��������?K�f��{���}�пYB��E��8|��tݎ��Lk�Kj'��X$�v�;�4��E�|PL��x��&�L�3O��y55��_Y�k]}!�l��Jm���ŅM�z��5FA MJ�X��� ��!EH��	��Oe�?����'��L�C̥��Q\�"��̋����K��@�r<C�M��r~:w��`	��#Dpd:�x�h���D��A�jAJ�H?�#l�V��]�-�]/�].&'�R&���U��e'��Z�̗>k?��_���m'2��dl�d��Q}�U�tޡ���%�^�����w�s8��c~/`�+ʫ��.d'؍���qk�B��,{5�Zߒ5"R�B����ŀ�z��B���7��uԒڄ�
�@��Em�*!P0��VZ_���u����喕sOD�t�*�Pf��E���977蓘X��@����\�22]�h�u��P��z���˔��!Qv��_?���uw)�1�:�ND#��
	��o�%R%P��R�_L����s/� |�PQ��GV�`KIQ%
�~���ib\{��ux�$3��JRd�LIઔ���6R�2�¬2iiٳ��٪ʪ��J��z[]_��o��V�'�Y)��:�'A"%��鰕���+{�#Yih9��/0�r�"�� �V�0E�C��1Doj�:6��Y��"��CГ^hՔp�!����7D�!���V�-	�:�����nQ�#R�V�����l���S#��l�-���$Qp���6p����̉01����c�< -'�J�+6!?kvv�C��h�؇���D?�����:k���߿�5�l���{4�_ãk"�/��%l��?I� �^^���!��_�ٍ+7������""����S=a��,���դk��!DD�����^�Q���Q��!�� �Ky��A����2��N:�M}��f�1B�m�l��ёq�����O� �	���g�8�5�u��i;{&D�g$.Բ:B�S7�X��c��u�|Y�CQ�B�!���'<��G4<t���!݇�#��|������,"�ζ�XU��4Jyuw��˟IXkS���?����}O`��9�r��"�&T�:��%�%ܩ*�MF�']���.և�^���*|[���{&�4#��LLJ���V7|��e	��Ԓ�c��	��/�kv���)`  {�DB`��䢸�'�,h�7ukj"� L) �#��(��Iue����`4E(1&BX&�639!bd��A"<�*�"����YCc��he�$&�+&�YP�BV��;]}=�w��V�>c��~ߧ*���JƤ,��y:A1�5��b�X�A}ܴ�jѸ!dm�i���>n��O������?!� 0�x	l��h$~"�s`H�K2`�3����0'֌����H�����kQ
�K�B?$�Pa\F����8�v���m��`�hK�s␓Uؼ�n� X�VJ�F��Pl\��Z+��ˡ���g�E	��K�VW�7��^�
^�6���jt�?�\�g���U2���x��ux��f6i�lo�O~"j���׾6n?�$(��{����$ ����'R���ڢ0���%K�R�e��=2Rm�OGD�S��	�*��""����M�#�𱌥�����,6t��FE�m�%d��MY"����:���Hð�qL����ΎF�w������5�FQQ�<�M�VG�����6�@n��k�u{�$d.ĕ��C���M���ҩ'Č8��!n�645��ԡri�Zki���k�/�W	G������VF�g%|�tr�B�Z;��!�[����g���W~����������7�H��i/p�������r��0���Ѭj.'f��;��Gh8�,����94�a}8"���%[YZ����s��	�#�L�Kx +�PQ������O��������1��P%dSo+���<�Q�X	?`�9F?�z�^ף���sK�V>7S2y��Q����X|QSʹ�7����,�v���B 1!d�1+�i.I�U�皛Bv�T���=���?�ڌm�-�[�N+w �H`�uO)D���g�f��-_X�"���?��O�M�g-*�N��-,/-@:I2�p�G�ϱ����V�£2�����&ԉ2k�cݚ����e���A<,˦�%;��H`+M�IC�bɈ�%�����6�`�"d�=����o���mbdA�5C`X��8� +)����b�������O%h���QUQ/b01{Ț��,�I=�G�Vw�?�`j>�_�/�__f���v��5�����L�ʶ��{����!ϴ +�n���_:k��sz/���YC���ޯ�m������w�na��'��ɣ�z�/���(ȼ��Y4�B@�b�a��PH~��L�G�UW�ř��E��'��$.���C��O=o�n��xƕ�)P:�@VS�Bш��!K/x�6��"6�}Ն�m�R���TȚ�a���h�޿쐽NV�<BBB�����kd�08|e�t�z�Y�	XvJ�c��&�}QG{�MO����!LXl��rD�v���<*�a �1��5�J!�$w���)֨������Q	/�H���#Ps\1�~��^�����y��UJ�ӟyyob,+�Xo��:��"�����'�_����Ղ�kS@I���dyJ�E�hs��3ӳ����dR#��jYC����|�GpqO0��Z��p<�>���E;��E����y{�[o����M�QgjCd�W��:B�`0���n�i������o|�����LΰF߲�.���nk�=h�O[,t��64�-���S�}��Ew���A��ޕ��=#��Q��Y��w��=)�!�,-�V)o����]�>n[�h��ُ��'iO^�qY��T����{��w������^{S>Ά8�%�9��O��E-^�Ƥ��t^���Ҥ���j�[�K�V����z`6�y�^�_]So�;k��w�{��r�Z�I9"da5A�b���l<=�XW&j�o�6x�+VUm\sE�\*sO�05o��oڃ�u�=	y��!�6�
x�ʠ��=�R	@!q��ǿ�9>���8c���ƈ~�9�a�PU���l�Y"��� J<,~��سd�d}�{�	��	��hP&!ӵP=��]���H�I�x�X!�>|�S���%k�ik��#�H���t5�X�\)G9��y�\^��AEX�&����3��oB�����y�0�@v�@�P�SV����m��9l�ϟ�W~�㌨�����:z�����}�^������~���x�f'��}s���K�D��>Q1l����sv����w��k��qeM�ں�����XcU��H��7Y��ݼ�O,Iة��&�lAT�'�!YX���ӭ��Yf�e�ڋH+^������u:$է��I3Shtl|N��kОG����>�;%�h]Qo�d���������U����A�-l����x���0��,�x��@Hό�x�_�c�I��y����T0�$������	I��^��Kr�5�bDы}��]�sG���Y�AY��Z��{�F�A��&Ȃ�Yjq�V���k��D���)����݄�	�욄T��k���~��s�[-$��ti����%���X��#Kb`v�\$"̋gA ,�D�o���ԔZ�~�CY�g��
���`�&)�iS�mwm�j���k4�I�9p���܋���O��h _|}��X�R���E�tŁ_%x�����%Մ�Z�h#N�go
���j	���Z��{���� �K%�^��ϼ���+�xy$�m��%���gN�s{ڎ��7��j����z��ma6c��k�i���>g�����v��H
�J)��7���G,�8o�?��#S�����ؓ�^�';-����b
������-ݖ�?��]x������S���Y��ѳ��o��;'�l�;-��C�����bj���-�VmW��F��Q�r�r��e��@*Q�57�ړO���>��n޸+��K�<*���r��O�u2vk-�	���+a6|G��yJ��Q�܇�Y��u	J���=A�{������[�ػo^���]:���)����I|0bCCl"2#�6c��9�7g��`����ؘ��OK����Y+S�e��������1�+:�'��h10�����{c��ZYQ��6�~b}��5j,��Þ��H����p\|,�uڨ�aAhVsQ�P�wcu�x�F���t��ԕX��W��'�MSPh(+���/>wV~x�����{6;�uK�8�Y���Tzu��e�D��[�nD�( ��+�1ag=lI��n�����4��$wmSfrÓ%Y��Rq&X�"�W5^�3�u:���`��#�ǩ�U��@���}�	_�O �K�n�Y]M�q�����g�Ys<e�h�E�:�q00ۈ��l9�n�������_!_����_�[�ɏ_�d,,��ʆ�M�Y�$��ME�v��A;v��t�!ww6mjrN�f������`��5�=\���Y����밈�\[��y�}�����+�DS�©�u껞���Oʞy�qkoO�����	:	���vG�]��>hs�����o�ѡ�>CO~��=��m0��}�s&v��ɛ�vv��i����~�^|�i;��1;z�?3`�?}��#'��̓G�}�1���O�����.)�f{��	{������ФE�!����r�h�Ũle���#�����5M|�^m'� ?�v��d�Y|����Q(v$D���&#|F��!���Xº�F��F�!p���3�{,��*H�'?KMh*o�R�L�WɛqI��J��~uMX��j���˙#O�L!c���]���jjˬ����"�MT��Y�������T�qig�˃	V~c�}�M�i��֊��cTf]�}�K��]�������Ϝ=y��sӋ��� ���B�(m��.bɨ[�����,b�rY�uY�¦5j��J�v�i *-�޾g�ݾ#?u�Br�Qc�F=�uA�BQY&+X�h�={v����ʂ��hwW�5K0��H�d��c��۩�dq۬��M,:���>������k6�p\֍$T'��w"��&�(��M�o�\��� B�y�a����{��rH��#$#{�ç9�uID�Ͼ�嗬%�����o�Q�`�Ɵ��	S�n���L��L��Ă|S���͌fU0��������ڗ�E;wZ�`�o������o�2�����
�ǲ��"P]�m��+��sg�������~;$ez�H�;~@�Q�ݻ3��oN)З���D � �?�74!��#QY���g�N�	k��d����v��a�uÓ���RNOm�����u�P�CE?pQ���QE�:�$��Af9o����ۑ#�����X���Y�I �s��g�&^	�2? L21ﵦ!@A��&x���w���13�^w�����	�Ɵ�!L[mO<u�FG�e��l��U7)	/��L��{˲�t��)���V�-�	���dcg�E��͵�uUDߖ��@�C;ጝ>����#�p4@k�.�������;�����׿&+t������.��CcV�-ۭ�����(K�[�9d��l|dVz�ܺ;��ҥ+�ppHL._M/�J�ҵ��ə`_@Ъ(&���o�uo���KN4?/�ĺ������a-x�3]�cB����v���9O����U[֘˃�F/Zk{XHdW��
.�<V�'�F,YgwR������	l�Hf�����������֔�V)���f��I�a��������V�Xu�E�
�K������{�����ho�vݣ��՚�OΌ.ۥ��Zy��gn2H�B��-9���������M���[�)	SX�t�n�L�O@��_����BQ�L �#\�2�Ý �Co="��x(]����&;V`>i R����#|@h��<nNu��q"����Q��' ���?�O��v,��@��o���-d��/����O��=�� �p�����f��r��["Z&KVf��vL���rK�X1�^Y]֒Q�ho�]Rr�Wɾ����O�����3+MfgǴ`B�&kD~_sK�Ν?a]�L����8(F���	��2���O6�'?�=�T���-���m����w5����wu��l~v�>|��-��E�p�V
8#b�h[�V�3�L��#p�� �p�)��c���F�p�1���9<!g]�2��3�����+.R�*���y:.�����W�li�����)K���<�����CHHep��l�X��s�*7�BwLO�u �X�Dz�5	mT��A�U�S����0&�S��B��#�	v�Ճ��c!&�'j�J~CȆ�*��Y!�h�!��X"@��Z4!��t�<��;ytq���!V��s"�Ը�����o��/m�������_ �\���^/���i�.�	v����Y,��	�<UdvrV�������b�@dov6#BI@$�t�9�X:!fߵ-YL���������K�.d��y�3�Cn������͏��7��mY��e݊�zL@�¡���6"r�g�ȢJY�s떜�k6xw���>�U�Z5B�v<�oM�V���u�pl�C̕�^�IS��Ŏd]�7TYCx�3?BFC�|����~������R���!��E"bڈzh8D'x�����#��3�bu�z3�E�(�<r�ͺ�h(�c���,�o~�����\�i+��E��F7���FHe���̞��"ER�"���ztݺ,��:��S������f.��I6�}j� �$ON��Y���i)&泲v�v�����-�h�Ce�>i�����/��kjn�n�zR�#���РГYܢ=���H���\`�BiA�N]O�b�	�p8���?�^�$�{�k�
��5�Y��tF���UiX�HvA�)e�U�[ޒ����M�Jb�¢-���Р���~�~�?�����~h�3A��PXu�ȊP�Y�5z�Vs*eebXQB�#k�|t	�J� ԛ�qq��^#����b�
�E�F�9;�ﶴ@q
�6����@j��'���UL+�"�ko��v6x��BZ���$�`i%v�D�8`��)�v�"]C��bY�,�ϙ���ļА7���PR"�4_��e?K��a�l��لp9'�~�9�)�vu|rt�a0A'���9"��5�z2��7	b1ID�E�A�>��Y߁��C�I1�L:�#W�� IA�L(�M�k����8��Ĥ6ꊿY�� �J�#zF�Μ鴶�-N-���I�smDp]����N�pue��R �Ɔn�/��ɵ�6==mw��I�~`W.ݴ���k�����]�~Gʚ��f���GG�3�H����4^���������+m�\���9�(E}�-�5ƒ),x�!���T��:W�@�L3�%�&Y��(dd(�C�5������[��'I ���Ѓ��Oz 4�ԉcn��ƪ�5�/��s65?i#�S��625��mZfaQX�(,�����kT�j==jI�mm����`q���s1Ni�\h���:^���b��+��IK�8s�٬/� +�i�	K]��+��]UYk�u1u�u��y��O^���s������v��3�x� p������ )���+����P��W�04��Ҵf��I�&c�f���EЪ,�ʺMO-H�(&�e���J:�p]H�e=��E��ְ�A���:�:��ј�>X�E�Ҙ�ɲ�/����}.���%����
�F���	�c��^��{a��_X$J���H$�(+�&�'m5�g��z�]J�eA�(��y(�J�{���v�֬�/J�KI��G�VXV���|����,ۃ���m���R��e$�(]���k����MI��5��3�43=/TrӮ�?����HX\L���K_����3+9�r�b�H�ȄqF|
]PN�a��\V�C�b3@����l}���� ��'��	�S	���O�֣}�M8�׀q3 Ѽ:��e�.�C
\!����PXsK����K���̊OG:QL2�Bs�Xb��U0;#�OCS�0j��tuٳϝ�{7�h�oy(�ɋg=��$��R@r�n��CǏم�ٱ�����v�v��1;���g�t֠��P����q}�N_8!g:�C�`LvLa�����Ò�=�~�Ymâ�U��!T��YY|i��c�@B 9�E[X(ɚ���D�?�m���-���K����ٕ˷�P�� o�z'XM��*�􏌄 �)��H׶��հ��h�}\K9��D���/,�����Z6��b1�FЫ��Ӟz������Y���'����J�A����]mJY$�c-�O����Q� n��-v�p�ڂ�Ը�
7������]�dxT|`�sj}U �����5j;�W�-O?����K��6�pLp^m��Z[���:W�?���֛@�m)�ڳ��Xc��B� �cѬ�wB�bȪ����` �FF �?���Q˖�P���u~aEww׫K�E�˞��IӼ�W���Q�w��$	�s� "��iA#��x�M,�XOFG`
,0�$��U���h��s��F"rSQ�`�==vQB6t�ݼr�#M�?{���$�L²(�*���U;��F��ueH�s�#\�s6�cc�������ư�\�C{���֞t�Dӹ���Y���n�!VeI�"hS�6:c�(X �!�5�xsڢ-b6�Ϛh�Br��1k��nK�����~;r��.���}t���pP�C�h�DĕR!OJ��@�h�VhF}�:S�3~��\���b�Rh���6��A8���O0�@�h��K7�؅'��\aww�9�gG���n&G��۹����������	}>y��:�k'O�CG{u�}>l)���=m�N�r-�Sg��Z$�ׯ��-C
*�eC[���x���oL� ]Â�'���~]� �.#�e�ں���dP���sl%d(l/��{`)%��ڲ@�X��Py�i�w�!���)����_�Aѐ�0,$tV��)�r�1�!��$`-���t��,!n T[�[l�MȒ� �{���5h0 adt�JZ�,��l)k<35�NcX����B��z)u�9�I�k.L��~%���XY����ڳϞ���v��}_�s�3���/��5�P��=1��glɇ��7޲o��wl���=�w����������#B��1�d����ܓg�q���B��&�gE����llDB~B�#lG��_��d��~�=�<����IE�ʂ>��9{���){�	1�9���ܹ#6 �(�_��=T�2�)� F���~h�|�H����R^$��,��^�P��"pX%Xg1���W)���1L��9Lv!�f�9>�4R��G�ք,��������qY�W���+w�"��a	I2b)фHJ
%�6�+NJV��)��ۯ_���#�ٞ�z�l�p��a���?��{��f�d�) ��n#��/�bi�²�����z����]����
��}�e�7�wlxxZ��ʈFu��X�?�نx��D.�<��!��@)|)(��	� &�ٗX�����,FI
F�q�[I�0>6	.���12�j��FR���f�B��g�uA}}ȣf�N��z(L��F����`gd�	��(�铝����_��0Z
#)�J�����e5�y�_Bv��Ō7�z����=kmM��n�?öB�wL����0��������a�i�";@�&IVK�6J��Q���w�.ɒ����&/�扰"6#/Kv���? �5�J9#f������ব��8��'����k�x�f��^�Z���E�7a�����	����η�k|�Wf/�E�%(�J�\ZR�=4rȕQH�~5�AD���`�Y�x�&��C�<�]�Gp�C��p8sC&栴w4Am�]�]���ݲ�^�>|�]y��|�a	u����1ݹ�X�*	����J^�H�"����ߕ�����O�i�53���Y���]{燗��Ñ �)�)J��&��:�V���,	���%��D�k��޻f7�B�{�Wi&ꇐ2n�;��%����-�O�q2��)����"Z}@X#F�G?W�.�,U� ���e%v�teP.�\����@����O}��{C#�*r9����|jQ�҅��|5�FG�(U�-|DE����kH.����&'��R�Q5R�ׄq��}������>n��e`��p�k���`�.|�������������ǿ�Mk�j���bgN�{%�K���߻j�,+�����3���M�n+K[��[_�� ǀ�uۃ�m����=yᐧ���Y�avnξ��w����1Y�:�f�-���>ͱ"���C�D�Էj�=D�A]u���E�PXE$��+kS%a�ֹҶl
A��k#ʒ�sK�u��̞�H(��2�P@��W���[���d�%�%>E�|!S��Xrf�E�Q�R�&�n4���@��`-���yR� �Jۃ��և7|��-��{��������|`����T+~�[��omF��Ǟ<�n�׾�5	l���ߘ��y:ї�>�
�I�����P |���:��v@�\4�T_�@��Mv�Ɋ���:�z���S&�%�o�G��0�§��c��X�����Jqv#E)N���@,I�Z�]&*�(���4���ů��j_E2�>	���`6�K��R*>��RN���Qug�'Ac�Ւp��/a��
�+�!���$����4)�8��v"T8��^A=��1@P����N�J����Y��GN�	����I;F�;(!�u���	e�9�޽!��g�1A�e��9�!K$X�)&(���ɴSǬ6�`����?��� @𿂄=#� /�PY���E�=4n#�H#:�fWZn��m��e7i�ZY�J1F���FJ�+�H���VW�N���Fe�s]��_���c�s�՚�"z3����'�㶊V�vO���ԙ)!���!����E�r*����,�R�,$�T)��2#q�ƋdZv���j���<<]3έ--B$	;x����}ў��{\�a�ś7niY;Vn����Sv��m���a�^��_��]��v�),�-f�%d�'���5z# �t���<�����y�_��z̵�Z���PL��9�n�s��:�{D��7���o,�:��0�)�qDX�AU<�`r����I��ź�=���3���$�//�d�Ȼ�BP?�қ>�W�_��ex�lx�����j�ǺEܤ5�E-.l+�p<��M;aO�ރ>����H[�\AP]&L�0��dW��3���{B����O�er��eE���i��q���ə)�'lva֦ey�Pt6�_��
�nJ�K��żL�o��c4�8y�ۙ��✽����Z��W��(-9��b�{bF��[}ܫ�3�X�U�'Vm��Zk�7�&�����%�/%�T�U�y��*��;����_�����'�K�{�?v��kȿܖ��a�^|�z���$eXUV/�=wZJd�&&K�h�cgOhܪm���D�<|H>L�44��4x�_{{ZCd�M��UkHd�v��L��8}����Y���:���;$�`�4�,-
�}�ʄ�lS}2����+��m[Z�����|�9)#���pF2�q!�3�G�t�+ajp0�H������ �k����>d	�W &٠�=a�9�B _"?\0;�q���t�
��'S�`���|��z�,arQ�R)�Z��d�|ڄ]��J�VԘ���<XƔ�����(�rw�$jy�dI�5�}��J����YRG�h��e�p��]����&@��QFAҚ�u���Rg\��L'�=�}��hU=���'�3?���⎩��%{ �X^_�
r��K"��eE+m�XA�dWױ	^>�"�� �}����zy��ߝ�E��B��l��D��={"�g�ԟ���gQZ7�'��A|�z�D����7A������j�3V~9/X�iq9��ݖ�i�Tg�%[S��u�CB&���ۚ�m�������Q�
F�y啂�є���'XD&A]M�ϳ]�����X�:��DO�]�,M�g>��u���9�h�Ξ>i�p\L"����5H9D$)�f!�h^���&�A�n���PF%�j@ߠ�X����ہ���9�ng�vYooJ̙���E�8D��Y�<���c���B;?꽍r/���!9(�1o����$��TRp4-8G� `@�)B�X?�'2_:j���^�h���.CpC8�B���Ů�p<.�@`�U(�TX�/�h�XZt�߬*�Yi7/"���B��4�Ҵ�����\+�U[�X�����ۣ668esSY�Q�ԹTf��zd�3��$���DD�,���)��@���A�|@dwN5��`[��lu�:��[Ĉ��e���|m��ج��F�7��z��FIβ���MO�3Y�g��z &�D	H�X�����J��޵F��Ji����U����m��s�S�|+i^2��əS?;�Z��@��?h���s������O����~�����W���_�_����Ϟ�ゅ{�)�����`c� ��&��P��rfъ�X����$
��|�Q\�P�F�M�R�7��QO#��b�m��b��O�������+����~��ɿ������O��W,��ڝ�S�����?{��쏿n����r����k���,��%��Jy���wFltx�W٣���v��kDĉ��xza���@������t�	�H�0��=��:�������r�R+�5D��\����q�;~h���=���_܏�v��T�b�P���3"ۥ�`0>�Ɔk�� ��/��O"S�x\x���	�D�Z�wj�C�u��Di�B.�-�Б�@]���v��A;u��oPG�,���Zd| _r��y�W��AKBD����\.�㄀����5�\�hMĶʪi;l&�bW.��շ'��(]Æ�,�	М�RX	,�g X,X&s���A{�w߰��&�	�������%�~ ��GT�y�]��xtt��+%�H��?D��q	�Ȝ͎e)6�������jU[�Vg��V�M�����Ͻd+�E���W< 4;���A�L����^��ݹ~ObE�W�C������.����[ұL6��0�r�֘=�Bi�S�&�.6tĚ�V�Y*�l��6�LtXS���ᴝ=q����;��e��?������M����bH��`����^nqٙ,����W��w��޹m���WVէyD_�a`�|������o�Yc^K���ŧ���3<�G"���K2�o���)��y@~1� E�{=ǡ��2<����B�s����:��8��@"��YO��D�+,$ӔJ���hH|�k�ξ�b�=�#����6�`g�Z	����<��`y�F]� �?}F~1���BǛZ��o�e]�`�ׁɽ������k��t� 2v86�b	��B�qV&�,��������C�#1{���v�x�����9����L�flI�UkK�����)+�4@�r�.o����j_\D�Z6���L���n{��uIVGꭴT�9�����;�Q��cō��^W��E_�B���z�U���/��Ko]�?��eo��^��{�m|l�F�'��ko����[�;�f%<wnݳ�)Y�)7lbl�ff�]�z8l7n�V_����>�ٹ�Ϲ�P�ڕ���&�����ИMN���mO�sc�.�{����{��W��nz*Xgw�ݹrˮ^�b�;y۫���>ō�[[��'O{Pcxhط��.-�bHHD�)�^��^~皑`� ��L�<�2�u��a\�F�/�bj'+����(����y�B/��%��w�����o{�EU-��R]���+��ҵ��e��dKܳ����x[	\��7[Gg�?�^�U�2:,&��1��	�cIk%�L���^0�Z0�a�9�(x�`8�QROĝ���M$)��R���%�b<	`Apjf"c33�6;?/�
��(ьCz\ =�@/���xab�W�tNG�|�#��hdE��}�Ͽc?��eiӢ�겁].��[��:�T�հȏ�W{���7��CL�.4�C�)�BZ� ��0ڪ��Y��I�D��eu_ I�)f�p�����׍���^�ڕ�dmI���e�f����y+�-IxVmbj���,��`���Ib ���e�F�Dj�ơ$���ܐ0�vd����*e�<�O�@�uU�_p�(޶ ]f1�>�w˷-��哕��!�)�(�<k��y[���N��ؐe�{�ܕ�w٦+I��s�4���z�$H&��x���M��sgO8�ƿ"��Yo��è�O��cA41@;�xxs��"`�`b���,���~��z���<q]�ވ�'��^܃g��ÛD
+������Q��2'����+�'%.!_<�1�7J(�f�%�mJ7��/m����?�� d��TȺh��5ʱN7�X2�$�F]����S.KG�렘��o��Q�}�����}�CdD�<VC3��|�?�j���i�����\X9\]]&�^���7�߶��I�wu�J�;r�׺�Ү!5�z8Wf-�I{���v��;z�K�"�������Nُ��ǭ�=m7�޵�>�c7o�_Hi�.�0����
�V�1��We�Z���56�c��_^.�,Ix�Ű;�)�!ܮO@%
�욬�J�0�,��V׫���y��Z��l�-{z� ��������(Cr/}�;�AS���g뿃#߲�N� 	 �tH 	�=ʻW�y��L��^rz�d'v)qW����x������pMhEr�����L�t�L�t?��U�+o���	 ���\�V�D�
�̟���c���s��_p��-��B��[,!
�-z��B{�gt	>;J��wg�}}/�3�uMd�)D��<�)8N�%Ȧ`�LL��Q�c�d"���g�s���~�vg�k�QT2[��~������~D2�E��(uL ,�C���H��gan���=)x��q\|*�P�'�Z�a��P"$�F���W�Сk�v8!X��@!H	9��bC͏R����;�E�%�䧉��X�m�r1-e	B���j�w�H�H۫�^�����0��)� O��[�(��2g����蒭�w<�J�՟�ۿ�_��mA�]�#@Н�]_ڱ�����ֳ���=��ܟ")�e1�n�������v�����o�{��m�Ȟ<��YjN�AR7{�mS����$*�˚l���`��AzZHqBl`x1�.��1�|�b�j���B`<(�B���:�>�\�PJ����|���w#��y\z�-��t���= ٘�	�%"���aa]��?��۸��ͶB�m�V�L����?ɹ꜄功�1�,��$}ǧV���yݳ �\b����/��˯x�"<F;$�fƳ���X'�v[�ph�����	x�";��y�zϋ��_���Q�$`;����4ŞɄ�Eرne$m�`���D�UW�}E�}�C�;>J��~+F���(N��T֪"���`U�`f}����mu�O�1�����l��2����=�*,��1�-�{C��h/���`U�)��uuU�
��Z5�( ڱLP6"�pI�ħ�����.�mz>'�c���}j�'<�_�{�6L�П/dyÖf6lu��t@_��v������o��c��_��ݺ9$_c���w}۞?_�gC��#�k�;�w�y�S� ��RZ�FKS�m�Erg\?�|�pg		c��8W�p�c�9�U�񗟃��\�j����?+<f`i�W��14v��y@�c�	��YG;��]�X�|oOL�.�*Amv������b����v�3�SS T�Z �Rk�~�˾�����7��x$�Y��2����[���������'?��]�vA
��2�����D�P��U*Y˲�Wڙ[�p���[O�@�A'�rp�Q>BY6^А�#u��Oݐ���.�n�k��`�q@V�5�Q�z�����޴7_?c��xM��xg� ���`]#]=���_�3�(�@^�+�Z�����	b��S�幅��40z(.f�d�4�?�'��2��vF_�X�p��)#G����(7G��":�����V��7^���O�\o�}����b="H{w����w�u����/�h�Owێ�ͣ{̜�KM2���@���t�&���|ͨI��_]� xY0�%�W��{�R��ԧ�h.X:yY�j��+Bn�H_<�H�)��565!|S�����.!��E�+�@�$���%>:°�Pq.�㟄��/�r���t8�s��	����������4�_����c�#W% o	���쑵�vڅKg��-Xwg�>wA���:���._���ݺ~�R<���'��/�i��3����u,�O+�E��������s���k���Z	���%�`�`/sj�V�I8Ϟ���:��W�g7�KhDo)$�F�wR8(E�nl}1��F��A��5�3��WW���'$h5����V��6"-+oƮH�����]�4r5�i�('�RD栦���B���faߪkb.I���>�R��_�jo�y�zz���6&|�.l�#�fr3Jy%��P��gE"K|i`�ݣJ2�hf���U���|b"ײ�]1D4���/XW[�t����3��p��/YC-��.Z[�%/Xc�Y+ީ��Vlϋmx�@���n����^�L{��]�aLm��w���h�Xy��ݢ�
�����:�!jt.e�eD"��Ή���?au5jG��rx�������X�{<w�����]��B#+%:��5�r`�p�>�	����~Q�
���?~�����z<�(� ����y�:K��e+�
(���=��`@aШ��}�-�����m~rA�0�Qfs�}A?�	�zU�a�n}|[��e�t�zϞ����\�Q�D�&t�crIj�3�c/-���g�⬾/���Z�`D�k�ς����ҫ쥷�ع��ڵ��V/�p��]��VŻ�IDY�]�Q��Ch� c�+�� ���,\��JSt��A����C��Z?�EK���N�����̬��j�
2@�@�����:���'!�S'����e$Ք�dm��dZ����$jV����	[�/�\��͎�e��!��Q}���^d2�����5�Ŝ�9�jP�Qge6����Q�jᨲ)�z��r+q|\i���>�e�}�I�=�Ub�D���=��ߟ���ϊl�YL찊��:�[YD�*r�J�NKWv��)�5A0���{���ܧ�|��j+-���ޫ����(�\� �_�x�i�3Vju�V^rբ�+:�[ߗ��`���?u�<�->$�
�����Џ�] �/D��!��;��������.��5z8�����ѾF̓d�Γj5M}�u�豁�^��`cC�P	32��Wf�Ҥ���%[�[��7��I�g�����^y�57���s�v�|X{F��x����.\=m�]-V.a��m�3:��&-����O�-)��!k��������Kvz`�+V����)�wK��p�����<�������"��B�9�AA����`P8DNu�H
��k1'��lM���/�^���_=����N~cGpL�,j Rj��,���N�YoW� �>��:��GwlnN�B\Gؓ�2(��*�2΂��E�\�GQHV��F'�bl.����^�I_Y����z���jl��	}Zc�S2��=�v�@I���S2�aj?�D���{&�w2���'�R���IN�9�a7�qN��L��h�����w�YL��;��_D���D��Z�ȗM\ �<z�"A6찲�~т����:G�8��_i�y�����?�)�O.�=ڛ����>��zAh�5���߰��{to�xPHN����S��hg���~$�bE���/l�z�Q�W_�(�X�;��ŅXB���3�.������%�+/�Z,��j�+/����&�{l�+���iu���E����Č�_ج�۵���Ĕ=�{7ۍO>�ٙ	���u�\KE���Et���e%�
|��dfH�h\c	����ƍ����*�Y�ƚ6SN�5>:gc�.\�a�/����=*+��v=Hi��|'��ɖØL��ُ���H�F��6���y�As3����mye]-&�F���bq9�j&�&NY� �(�]ؒPR���'����1a�:i]Ԡ���h�!;��	���u�,�)D0��*���;A\�0{�3�P	*Q2� �`.��� ��Vה�I�$h8���LFD,��Ԙ�0Ð���hT�´�0�����;!����(O��	(-?1����E�+�FD�-���Y� 0�ױ�y�[x~���'���=��Nc���g�\�s9�;����/��g�r3��X�Dv�.c����uu�X{_�������T�贳gz���Yj���m�k�=P��ް�����]�y��ݻ�Ć�i������.]:����$n�wj+䧉�l<�x��7(y��߳6��?z@����|h�VV�D��bE/H�c����(�`�X�U]S����qg?�R�?����8>�1C��9�"���B_ٍ�K�+pʕM�1 �N�dk�-cO�T"� �`6�.x����i�+����ؽ��ѓg�#bx�#9��b���/����dTQ�^b/*�� d�/�I�J�3sIh��a�K�7X}�_�����jVp�NR����L�]�Zj_�z��x��MD��۷te�N[k�IK[���$�V�6�4cT����Z���٬�����
%"H�L8^�Tۛ��K�0�v-b�)��+l���ޕ�v�B��x��^}=*�+���
���.�oO���&� ���y��Q
���-�`��[!�%�B�� [��2��˱n��1B�Eh�r|tʦ�k��L��~����WP��^����4K�j�NG[]��75Y������%�}뮭�-9�ʽ������Ȱ~?���i���t��]B{�܀+����P1L�p�#��f�ӏnx)>��:�4�;���m8�v�C%f}t��]����+&}�բPPUM��(�\�]=�Z7�~hK��}�'��!��5�Т7�l.�8�D@b�A�C<����j����$T�]ϯ������3�6%�<~��F�����l��?�C��&� ��.<���,IV1���1���F&�LA����nc�,k��V���{uN��D8�p��Ꮲ0i<���'��M����2�/�O	i�;��^z��^����6��������O���[��ڛ�������2��O�XR��o�?��#VU�,��/ʻ��90ơ�.j��{���bB^�T��"�[[۷�`U����=��� �P 煹1N�Pi�ZA	��H���0<c�+�6���7q&�����AJ\�Ys�"�/s�G�V'8�����������n~��`�#���C���G6<<%����Ƨ��n�O�m�`K��.+e��e�Q�r�/{�\� d����	j��4ipE�lݮt�#��̤;����Z��H�ʒ9D����#��ްF/��8��a~�s�[�<.�Š�,��կ��y�hF��3�P����}�U��̗R�#������R�M"Vk_V�d|.r�rE5�A�}�o�;����c��j��m�d��p���%�hL�` f�>��MѸ.�:?ZQ�BUi���"A���c��4/i�|�*Y��~3j���?޶?��}��W{������F
�KXJ��h�����L1�ɧ�|��>����'���n���?oۯ~�g�OC�wF�l�J�����s�c'��|h]dO��O)�_���?;���ߓ�eW�2-Rlw��	YP������k[��E/X����S\�C�<0��
=��8����[�9��e��Bu,�b11�&6�I�&�쭯]��WN8����1q���X�I)��S}�����d��O�Zω11�,���^��g���2��LG����7{� Yt������Y��N�N���QY�G^ƛ�B�ƽ��.���iA?�m��J��#�=�ć�y<�zҀ�	)p�$��l��?�=I�C�Xq@��o��į\���|voQ�$��y!�����@
R<_�
6�}�XR=22�9��)B˒�5݀ʺ@����ШCJ5��{<�~�Al.�+���y4����"$�@>�;��[wrf8(���i��N��o���D(�BcC��9_l�n����BdgSVei,k�	myy����}	�~�8#�/g����������,�V,KG_�z�$�����c�K�<��w�ldx�.].�r����M����,�*l	�7E/i�~��Εe��S_���t�`�u `0t�'|�õ�B�ݑd�S	PFh�\@>�Ǌ]�:����2������b0~�[�d��~fQ��V$Fdb���UZ�ŹY�a4&T��B����v 0�!顨D�Y4!˄��_�����?�+���������o������������'����>�ͭ=E�� �NJ^�9"�����?��~����`�����fo�D�;�pk��B!�+!�ʜ�|���`+�K^ �F�ʦoEA[�{n��?����R���.�빜�y�ì�dUjH�WCA&�ZGH��PgIFEè���OsO�a]�ˡD��h�$�o����30\�F$�Y��>t���̪�4�@�{�tOf��!�8}�p0 ~��i.j�l{;�Y��Y�sѤ�@r��I�W^�Edk��!|�&�`#���b��0�D�6��ղg/\-�t����c��EFm�F��ߴEgZYр�h�@9C0`�� E�"A#u�����l��/���/���u?H�P����@����)����+��:H��6(�x<a%�Ҋv�lrǂT槫3�V]S���[KsZ�(s+B�|�����
$d5��U$�]y1>(��MLL꘰��i��?���!���$%�X��i�G� ���u?�~ "���;/���wz���#�g-O�����	pee(&KFߗ
e�(s�X�*U���W�(0K�<*�� k	���.�H�8	..aI���I@�(�M��-�D ;j�C���d"VYf5u)�Y,m� �����ΉO���P�2���/F���j�k�H�hS�C�r��$I��Y*]Z�p�#H��Veq��Pc$,�ӵ"(�H�ni-��̡|)�Fb["Pj�'�2 �����"T��r2Ul�z�VA�FJ��#�}��C����K��聽p-b��v�n|,��	�נr���"heV��[���cHH��rq&���Q����G��y	%Q��X5�6��FO�_����i{6�̖W�̇haxVSv���$.xE0����j+S��h�+;�"�D��J�}���6p����l`��z�z����R�Z�"܍B.+#!!��SC���["�=:����N�>��]��o���^A�N�lo�����nu�P�NԈ��L�����*Wǭ��)A����#�ߌB���-ʭ����Bu}ڒ��/����}C�t�:�S����ưa!gr�@�nm
{J�nR�J�!��I���!HI��K��M�(g`����[u��,"��H�AGiV��h:|?�p8pn�<�'��䔓��D۔E��z���A�}��q;w1�(\�ٷ�{��%:���b��/�n���v� �9��Q���CXO��B`]�O��-r���)S�%���q�s{��䏷�W� �o�t��+���b!vn���i�߄��R�^���k,h���w�Ej/c�s�:��s�Or�B���ųv�L�U��|#F��U���Ծd������'���~j������������(����ܛ�CL���f-��ih�VY���ںۭg��ZZ�a	���FU4�-֫"�����ok���Z)ل��5ʚu�ؕς_��(%4"ʏ���x-C�5����R�ڨ���)�B��m	>B���|�_��ᢔ��%��]�U$�)VL��%J�tw�����.�&�U��I�q9�id6I��� p�[Y���|�"�%��T-"�����a�!Î ��1�)��a�X��	|���S���߉YE�u��r��Bd���<�i�O�+�`����,�v��E쫿�W^a��X��54�՗J���r{�Ri�ڱ���M9�ζ.TA!��=W*Tl��[��?Jvhg�(1{�W�+�u�a�ήb;}&jׯ���4I�1�x�̾��{�d����#������ z	^��Ya�}�<��@�}�����}���z��{�q��(����_�=�n,P��o�-;{�����66:g�K��_/h��/ a����Dm����m|d�����e7|���
8���Rl��f']��_~����O���/ە��u�^}岽��v���н�"�A4��w�$�N� �۩sg���߷��ƛ��+�쵗��b��zYן�ƺ�}��]]�.�έ���/(="�#��7����9��'�����q�9C6�� �K��劸�<!Weͣɬ`a����AAkLF�ŤC�L&� ��ƐI�u��e�i�r�8��`ʬQEhE��
�傋�b��GZ�p��03c�&��>�bu��!�Ed���>/���Pj��h$�@D1klB�������f�k"�>!J�= R�ٿ���_�ڿ�g����˂���#9�6	o��ĉ�Y�ܡ`���i�ʪ�Ӊ@B�ֹc/�n68�g�G;(�{�{3����?�?}o?DM�_�)9�>s��s�v���?�<B�>p8t�.U�t~P$��hw�����Rrl2�ѯ�����ĚP��Hq\��b��oA{����K�\������m+��KU�%"Q�����@3�8ɔզ+�]����u��{��0����KYV��l!$:����!HUq�}Q1�u++��b�r���u	VJ�`$Q �2Z�t��oH�`�(�W�b��ԑd�݌�J������oe��؞8]�Qⶱ�i33�khKk�56��8���s�i�`�R&���ғ�LJ�~�0w��v5aI U{��`�(A*/a����;{[^���N'�c��`�@��~` އ%��w�J"8�rv �zZ�N�9��v>U߉GO�3�N�4x�a��I�ȵ� >��Q-��z�Nm��t��"�T{t�ݝb��1��X�0h=�%f��)�1�|���/�:���yAt��g��G�h��0}8`S2Cve�Fuo&N� h�P*�z�S�?��-��Ѕ�[W����ҵ@B��X;�0��:���O[YX�~}�����n�~��"A��C���Շ})�
1RBV�^W1^\��D����!&c~JQ��#SL���O��7+,.��u	��<���o���Md��Aj��+y����V~].����-,��A���/���I�A� �:ݯc�=�� ��U$?0^��< B�������Ԓ��u�wZmS��j�GĶ��/�����5�˫�ӎ�t�[GJ��PuLϤå���k��K{I�<�gݽ-�`UV[�R�\�1.�Vm�L�edҫ�+��8ŤT�CC������� h����� p�G��E!�:��e	��3�����*�9Y�[7v��؋/E-�fgIVc��x�3�����[����M�2p����f�%	L2�A�_��(��Hy5B�%6<�E<���a�KW�]�Tj�Ev�SA�"9�E6p2"l~�ם<�l��ZZ"��H�$X�J^`�-�+!v��v�>�B�W�Dh�wJH��:�rF�
�AO�(0�e��܉x/Z�d��qgw�u��Yc��x��Ǭ��N�D�Z;!�#imY�Jg�ʰTp�T����9��E���Ʈ3+ٜmI
1��\���=�ܞ=zb��jA�G��@!P�� 
J��<�C�� vY
}hhȞ=y&~�@�0*9�E��� �7�(�d��i������T����y!��`2svx�tY�Nѧ���[[VD�ckS�%v�
m�#!�X��[$G���'Y�t�"��]��r��*�������I��-h��G�Ҡ��V�Ce�:	&�.(�H��q&�P����9/:� �ò��4���/���#<��~aY�Y�������r������L-���"{Q~عQ;y6�iQ##���q������ۃ��63�/G�Q����	�Ж�R��\�P�])�";q�TBT&�Wl��0A���}{��x9*�����������l��v��S���Xj/�,���._+��*��e�EG/���9�m{�1�G��@w)����ק�\tt=BuD��P�Y�	}e������s] �K-���f���l�m��~���wmy5�1!��x%���Ӿ��gc�*���v�;�j��T)������x>吩�.m�j1^cއ��+��6�|L~�cY�1���Ҙ�(/�&Y���� ��������o��䒍�N�z-�����TJp�� ��f�F4x����@8��8�M��0��..[�M������j��m�iJ$���iH��w��XZ��@4.��%T��=��@��������Ŕ�r�҂�a�tTR����2����9���ɢ��
�
7I�gW<�����b��pAւ�t�:E����F$�N���]� ���f�,��%bg�YL.Z�I����t��܁�i�F���H�*�������#sŶ0�m��,��s�vF�Ίmh7�����[�ч���{f�iwn����b��{r�u�$�K�F��_o���&�b�O�?�`_���>�h�>�h�>|ˮ�k����v�=z�����������Ϝ3��a��F�c��� ��}�3�Z.x�#�0 +�������s���Ϗ��*���ط�����=1�:U��P���v�ŋ�)��Ȥ5������'B�Sp�j�65<���{_��T���9�ȭz�����>�
��RW��x`,��9�3K=���n{|�n||�FGF|����y).Y��5������!�oOB�<�["+V?Еy;�c*���C���g3�=�k\S�q�c)ׄ�T"�U����C�xE�\T��EHj.��`�]F����ɯ�XkG��_\fY�4U#6&A��%ǳ,Je�� tO6��Q!�7b��3����{�c��4���Yp7���$�E,A4Gee��y���i���I;�:á��X��l�-��8g�=�{w[��\P���a�{r~5x��h;_�-a��d�/.���Ҕ�0E�0+�Y���x?4@��ꚠ�0ϒe�`��ȗ�qw����y�g~�Rm�$_��|.0�K��/�����/m��#	�qn��#����3���:H�k�=z��>�@'���	/��	!�H���o�r���@>�[𮭭ۚ���ȩ�5����Kg��&�FDciDJqO�&+������d��;��v��%|>8a�O�H����=�`-���,����f�+5X_Hi[eUBGچ��n�{B�&�ū;�N-��'aS��`��������F�H���O[����Oy���[�������ӱ��o�C��R,>�բ�:2�B"'�=�s���"�76�	���<<Lנ�!�6�̆rj¼�1�}�X_�o#�����I��$t��O�l�h�PĠ����^Q�],F���[b�)+/�p��>"����oQ����[�G��"��k1l��c�Q�P�yD���~y�(�@,�8>�Z! �Չ�y�9T%��@�P��ֳ�b��M�Ë��K�>�����y�E��xy��lo�����p/Mh=�A��ZxVx&����0��_�����zm���?�=�!p��z>�)����jW�]�Y���#�7�du�V&-^\��2khi���v{tk'a�#_|(߷Ʈ\��L­��'�^�v���̊�1�J�3�"(LF��	�E��+�x�N���۬�g]c�ZU�=������=$��z��9^"��"L���7��8bWXR��#�qY'�.,�&�i��c��6Z�\�!LEɒJ�H�gΗ{���*r����eO��De�,Š�W%*b2�,L��ӛ��I,['9ԃq�y��e4�=jа�t�5ԙ4���P�#bu��A[����}pS���3g	�?܃7bFg,H,B��.���'��_�"t�������r�5H�H�F&�#�4����PrH� dx�U�@�8�s&ڧr.?LC����/m}�?�d�%�.�j��F�eI�t�/�<�ޫ]�;����/�`*���<:�y'
�xV��z/��4��/��׿z�wH!ЕL��7=0������ho��^�T������+A�H�O�3i\X����%�͏�	VB'�K��M֫�+-&�@9��!<������*D�-�y�&y�9,�0D�]V�eE�nQpQ�x��~Jw��D�c�VU����J<�G]�=�ָ��p)�X`���V�s0�\��G��G详B<B����u�Δ�@�sM�������-�,-�e�+�V4(�Bq �D���BhB��V�2�$j����25��e`u��:�"MuJ��|4�⢼��he,%�#�݅��SV�!�;YS���X
��
R��CYR�;X
CD��Ķ��8��R�2�F�w�⾌d��s-(�<O���`�ChBgC����4A!ɒ�U(���y�XT�$�u[�c+쾧O���[`�h�����L��*��L��xai=���喝K��G�tk�'�6^�z���m��6�$��1²$����E!����y�s���
�Lϯ}�oh�~�]�`��NB#�giApR>���ݿ7d�}斻�U�&}L�B{��,xG����Յ��b�?��w����	��Ŝ�0������n�y� �	��U'�V�0���)6SG���9��>��X��W���'a�����K}��˧=�P� @���0�s|c�u+YC�X����ù����H;��}�b�0Y�n$���:aSҐX�d��mv�]#����� �O$FD�M����_�G�,��E�Mv���i��lhl� ���b�z�0���:E�90��n�U��˯�`���vKM����� =�t-̗��+��ǭ��ٶ�����F�T2�y@���ɱqyny�씉#�TH\�XB)4)6�c�����fr���0�m�hյ(��Ҡ#a�\`��~&�d!�bA����y�)}����b�p�����|�9��%�������U�NW��Ң�˜�.-��D,�ϒ�����`��Hc�+�m�b	�x~���Q�U�J�m����olyy���I+̋ɲ�V�j��s.�D��I���x%@x�f9h��˵�	���g���Z�ҕ)+/Q�MҋK���J�A�FP�Tc�~�,%(R[^Qf+��B:"w�|+��[:Zu]�-.�.Scq�h{[{�����޺d/\��`�NI��������ϋ��,����N^&���}͗|�K��*�1���^o]���ڶ�����b��=�j�N�C&i�+�EV�����
������)�֠��^�A�����}�������}X1-!6�n-��Nh��ծQ�="f�<ٸմ���_m�dzΞ���� qX������m��ö�tߖ����g6;����J�-�>��'R(Ol~���I�3��C�TZ���V��O��o���cA�);(���䊬��������'j�k�v��BӢ�J��h�9�0��a��VU=����f� �"�n��/�+܇�@!�zD&յ�R���s`x��BC��$X�����=+hl@h�}�dM�^����
F��t�b &.�Z2�v��a��O��F!T7%��+��*f�hE��9H�_��y2��	P�,\�S��uG@5��������K61<-h�u�Dʞ�����@)Ee��AM��ӳY!]X��ß]���#^��g(W\jk[�::�d���ö�7u�� |�%GyE_����s��%�V�l,U�*+cf���|�5�Ťm
2����S�s��/y��xShR��m�,�L���+�A(T�G��2���S/��	4�����r��ͯ��[j�6!����;�L��6��]Ցc�
��J��Pd�gN۷��7��`���_�/v��#;T[_����[W�^�l�P;��g7L����W����d+O�yR5��8�%^����7�o�+��94�W�����W/�VU����Z��w�y��6H/&��i;��XP�u��A/�xt���y��A���4��ƈ��l^�w�AC������L��KV�"��Boo���glazŞ=����Y�,(�x<c�^�f�������޿���ªS	K�%�@����O����%����m|b��i��D�������j��%�@���49l��.8Gq�s��^nP��$�2����b���j��~j�o<��.�D	�~R4��8�&�t��C��(���dMM�ND�'�uSS��Cy���̺���y;y�G�5cc��v���k/A`�zn����E���x� Ǒ���`H�Kt�$�f�s� s"-BM�[�����Y�A9|:?"8�P3A���¥�^lz���ku�E��@�űgs;�߇<D�<8!g֊�v��)AM�� �+�i����ץ��Jk����2��55dlbp�7NOW��7~�{�WmG>���9i�5[a���/V7s"����=1<i��s�</x<��dm3�+��Y_�e��޺/-&�*���$);w�ʋvB�Kmu�}rV*���q<���\�y������8�_��ϕ��|-���$X0���Z ,�>�[+*�-��uѧ�D�-/��гi�-1ᾄg�Z)-v���<o��Y�A�5�W[GW�ҩR�ﲈ��LJ�7"�S0\>/�u������_�Am��^ �	�-���n�u���^R�(hɡu�w��Ф|�y���!�%�;�]M��a���� %�c~w�µ�7>!���U�nI)/�A8��DF��ۂx�J;��N`�'3��twu��>�����BHے ���)Z�ɓa{�ݛ����#�� D�$*I���h���}��p0��(�A�I�q(�͒���g�0�3P����ӖH�g'���ޗN�>j� 8�00[�����PS[��<���5)�*���K�K�'�3��߳�'����56��]��k7�߳�޶�Q�e%�s6�tĦ&lq)o]���YV��ǷlA>��|<�DKS67�f��?�۟=���Y1����u����H�~G<����3�Ϲ�D�`,>r��9��a��ǭ������܍{�� �v�F�7J�M��X�j_	�m�m(/�[Kg�������VZ.�D�YQv���Z���z:,d�ኘ��{aT�0�W^j��7ʆ~���w�M߂u�����&���H����Q�?��^pdRZ��!�\����!���{�D&w��!��a`�Ó���uY!d*�ܲ�	���<��)#-���o�~�����HD���)m4f�����O�4�����'��\î����|�ʵ �@8S�S��`��rP��!���V�k���sy���C���׿h�����ɩ��-Y���]���a)Y���u��������7hFB�D}��\][Q7�Ț�<�bg����@pvʞ?�ѱ����b��ejˤ�c��"���ry�GBt;xp����c��ۍ���c	fA
 �G����\>���B� ����	��2g��:�����H�e�\��!��.Ÿ�N�5�=�8�ϥA:t>)q�����6���M�sc���<�t��f'����g6;%k��z�cs{�eZ+m�7�/s�f�d!"�C�.��h�6�x��:�
����d�����xkE��#��ku�ڗ_b��e����T ����b��'�'	�P>N_{�磠pI�����`QB��B��d2$$ԳhX	�d�@�e>�}g�N+x 5����1�!$���Ν��W�w�D�0+�ZGm�_S.x承T� W��2�|�AG�r�����(X0~� XQ��oK�p�ш�,nZ*Qc�R�}�g��n��u�w�ǺNvZ{�;�k,��"K�Ė��0���qV��%�EV�X-��T��[9�9(��G�-�@4�@}��/��N��T� �A�C�I�mj���]6p���p8�j+���fВ�r�FB Q
{(�!Ћqҽ|��� �w��ֿsAhl�G(���L#2z�^�Z)GY����譗/^m���XJ Lm�bX�uޕ�����-�deI��,��� ?�� ���H�gW�f�<�"O!�ϒg�{�P�G����� �r6]�A���sË�%�bϥ��sto�	�����8��[('��)��w�{P4d�2~�'a�b�A�;�tAiM�g�����2B�4����P
��%*{H!�H/��
b��lN�Q"g1�8�%.�|���/�X�-.X����`�1�&�s��h�xs�͘������y��\��A�y����S)9���q��K'��t��u���G��2P��H�S �̮m
�L��籦��{�W��.B��E��bd�?N*�;$�QDf_r���;�f����k������5��M�h�<�r�3`=π�>����7/��!N
[��{x1��PH���~?�G��o|f�L�!	��6p?��^뷿ho~��ԧ�ȯH�|���oB�SR���ԅ}[�Y���>�wv�~����	��@d��HJ8���Nt� _�F�B;:�Xn��X�E���(`���}�AJC�������TӵUB7��묨>R4z�?�	�Ɓ|Y���ª�¼�lP
���{�V-4��I_�ټg$��	h�e]�pdx �|�O���O��!I���(j)a��
l���!;�����n�QЄ�}�WR��cI@�H��)��a��_*����������Z'���ݴ��%+*;�V�Ś����k�������K;0�P3���P�yt���OIi\B�����?�i�L�����`���Ɓ�,o��;�v�S�n3��k""VE�Kp+��|d`�~o�Ć-ا<���F��~��[+���$�38���3P�����=S�H@�}�K'8�|:qY�2�8��C*� ���/�Pf0$��
뇶��TJR}��T�D`��G�zuuř���F�":6�$��܂�ٚ��X��Q�aKך/fL
V�^h|xa%N2/KY�!�(� ��G�|�j���u���u_�{P:��(��Zc���7AM���~�[}@9��D+�;΋���4��/.nrSirzYZ������U[�_������^d��yV	�O��,Ѯ����+œ��6�[2�d7�.M˻���U�RS�H�A�209� "2bdx�u,�g:����\�̙HpH3�`�!��@ᧄ��='�[i���4��͌/��ϑ؛��ٜ-��mvl�F�mxh���y'�-��+o^����g1�Ɩ�$��C9񲔇%�ʤ,]���ڌ d��lO��A�bY�Z���v؅s=����F݋0�l(���ڽ[���G���Q��TxB{n#/8@g[)م܃ x������(��`��@�W���3�������/ܯ����I!�gmn�h�F�C�Q�N��e�b���F{��+ƞ�����e]c�'�Uې�/}�5+ս�L�-�����+�ܦ���J���aH�:ꬦ�Z�3�m�d]Yf)ʾ[AOY|W�mf��N�Ki>���E��c�J��S	"�<KjV����u�%e��đ״#��ea��R^趲�j{j7e�II?�"xC��t���o[�@2��eW	�W>�!��J���JOV��sk%�I98,�0�~���5͖3B�L/�}�Y g�b�"P�s��^>`�$�C|A{�S*�zL�9S��;ҹ�$%!yI�&���u���́��Uu���Hv��B6�`bY��^�hg������~�p鄝�0`���ً�^��ߺj��y�^y��]{�]{�]�v�.]9i^8iW����g�,�{?}2l7o��@ʱ�D�@���%�
R�j�^������Ƒ_����xJ���X=�ٕ�kU)'1
t@X~��c��5��p�K��=����:��oD#)�T�hMV�ňz�*@�%�p���^z��o��˟�Z�s��lJ����ܦ{Fl�頄J�P�mh�����C������ȓ�Ղ{������bo~�%;}�_�/��(d�#�ٱ����K���W߸f�=����)�i����ʅX�VZV$��������h+%�P����G��b�Y)�R&�u"���� 1��妔��xb��@u`,"�ݝ�dE0)ETy��$�����KD@�w!�$��R�|.����5�{��/�K��f�+�?>`�8"�0D&&(CY9,%BS�k�w��!��|���*�H')\"�y��F=:�]˹�
�-�Y\��!�2+�hq��K����F�|���i:)���R}V*��0�P8詬駟ޱ��1��	��jl���!O؛_}E�t��q9vu�t�7�,.���ҩ���86t�/�$P	Z���'8���3��t�Ep���s�WG�kRb�޳�>~#B��a7��y����ޮ�xI!g�?�!���:������k,]�����B+SS4�r}K��%!c:hrtV�_a	5|Q����t5�Q��̯�l����1�_�AaG4�U���-�^s���M���e���ާ�m|dL��@�]��+�g����y����c�qS�����5e�m�;�$/D����̯q�VQ��:���BFJ�˯�v8���/*eٶKRd,�[���w�ޣ�!���@;Ԡy����d#J����j��1�9��!D���|� CG�ЮL�un�X�QP�Z�t"�{�K�XR�F�dV�f�ox>SD�d,�"ђ����SM����ܣIԠ(�⼒�+� �E�A�E���#q�~�N�����J��Y�|V��dZ_ϻ��WZm}�����ɽ���?�@*�,����7�_�nT�[o}��X~�p�A8K}�}+h�P 6��N���q����:�{q�[4�4RZn����Wl��s{_m�*��ybl�cU5�Bg��������/�{kh�ڋ_8�<�j�v���!�=�e��w��F�#u�����_��|�y���m�[\co���V����f���ˮl���y�K�x��*����,
?rA�m��/|�m���p��ƺ[]����/�����/��,Y�hgne�|Mq#ʣ�ρ@y��9sm�12��ʌ��,�
&��e�Ȍi�h�G���)_��{A��65����f��"��킋�Pf���/�:L,"�U�����Q1i�
�\H�b��--
s;���˃Hfp����o1�#�C���X7��!B��׸b<�#�]D�XB���ή޳�G����δ`�.w( ����w�r��s�p:�K6� m��(�X�م)[\�/�����I[X�L���²m�dmie���'l-�h���L�PJym�����J��������g,��d���tn�`>�O�1�;~�VM�wC�Hn��o� ��h���#h@}|n����V��h[P?���.4�dݟi����V+��)Sߚ�(-Q�A��<��[]c��,�d�}뾆y_V�H�mCV~]�;�[߉N���X�XMc�Z;[�e�̖�Z;q���$�d�Gc6�dL��صW/Y��
9]��^:g����"����,VQj�����,S�l%BPEI[�۰��9�w�mlgEf)[�,�o�B�_}'��b���|�ѳm	�#����Eh��9���iؓ����۹*&ɜ�6��H�&h���#-m��s��v�T����	��DbX~�e[��E���Ϧ �Qc�&�p��50��`$������<X��w��g�kW�4��1���ur��g"pD��G2��y�,��HI!�^LEDE� 4B�QC���H�K�e]#����Xm�� �ed����E�{�zv����VP��_��[��pKְ�W�R���۶de�^�o�8;�78�._0����a%$X�@U� ��\A7��y0-���������܃?���(N��u����bx��AY�I���)Y�A)�5��O�ωN�VY��	��|����u�p �ܞ���ż����gwG��nZ[ܑϴjsk6�h��}fc�����j�/��oVI$��g�,KL��@6�؜�	N�f�W��{�ɯ����a�����亭II�'JD;�Q�@�R�7�-����_�yX������H7<�#��!\��VX���Y��GCQ��F���sAm�+��HhƐh��.ʒ�G
i5��fΧ�^[>O*EfuT0����S�iY{���E��HnȀ���_Dp�@x�h:��Dga]��	>#G�q��U��&ف^�����d��1�zL
Ӌq	�8�� Ø�Q%;dL���0y *e��$�a�0ѫ�)o���id�aT���}�A��Xk��!0U�S��N��r6<2��`>�l��Xc/�pd��>����9Jhґ��O�?�J���,��60;��K����U.��^�~�R�K���Ӫ�R�Wm�m�<�*h6����<![���p����lW_�仗����\�
�k˰8\��9��΋[�,��[����g6:<c�9{�dĮ�ꆽ+(z���%�85>�n�n���O�@@E��	%(��/)�۟<��c���o �"���8#>`���;�b�DǗ���L�;�A}�_��"zI;|�J��{�h���e$-���q$� �E���}	
���Y�斶w6יk�5�_]C��z���
*HK��������<=&�*$|�E+0�<�,v2*c��p - C��p��m�V!�NCx�o� Q���5�7�L�Uu}T~��/'�}O?t��`@$����t� �E�qx,�̷6�#@�cXEW:ס��E'3�K�N�X�mu����C���%������I�X}{����5	�{-DE��Smb�:���N����o}Ϣ �w�l�e����E)�����MR+�
e�����SB��佸���N8�_�Yq8{��v�����
Rim�w�G�Lcڪ�S�H}:f����#�ejg�� d��8�/��H�'ޔ����;�mE�x")]c�=�驹�Ld�w�
BH벌��-������#�z��	�������Ȼ��m�I��n|���$Hy�ck�+�}_�m��5��И�l�4D���<;G<Ĵ�����ܜ���{ɓ����ۡ�G�Wצ}K(6�D�21U�JZ��x	��׾�JQ'G�[���	 �Qi���*k�\����X�MYQ
[�2 5�Ei91��0�G��p�uM��4�7ҘT��5.����1�"̊Vf�!U��`,+/�Y��⚩���L��c��~���*� �1B�&]O�	�v�~���`�޴�c
�v���t��a��3Z���Ah3
�L�#���l ���zf��9S��6�|BSj쵷/Z�V9�+�8���s}���^���m����|���U$Rv�s��^'ȵ(�V�S����Z���9��~�{o�ڱ��I_+��o�(���y"g�,�R/�iq!"rZQ�Dy�Q�![YK!�4�;�=+����i���R��t5�f�m]�>5�U�������J��V�Vm���s�ݏ�L�VVW54�A���""�zO���J9M1���ũ��Z�_��?�����T�1vXv�����
���x�q�၌�O!�	����z #,A�#t(M�8EcK�'�#�%�����D�	"`<+��O)96�`�6�*"���X>�Z�t�Қ[BA�r]�D�|&���Y���!��|���*j��O�t�d� "�/�������1��Ɯ��h!|���@�	O�������������+��kW��Sv��ikio�n�Xb��.�7����c���zx����V�����>>�Mv����b��0|G�o��)q����f�����v�N��'��a�n�Û���gO�ƌ�ȉV��Z���@���Y)��s^FmqjѦ�����Z{�\�Όc�ʭk����(��6���K�R���$'-Fn�i���%[2J�u�������Ǯ�kazٞ��g�Fm�餷��g�my~A� E�HI��p�~����<9���Ҥ�`!�"�
�>�z��RJ��簃�+m	]Mu��46ۉ��fW_ɖ��}����,�p�nfV~���>#��h�O�巍����mbb��,�����>�2U����0�`��
#� �r�AE<�`�x�&b,A]d�a�	��/���$,�E�$DM��r��R���#k$i��zgs��HR}]�"b0����'�F���-H��D�G9-\+J~!hh�Ri�-�U̚�$KA�����:���ڃ�c_&�v�3NK%sb^�Z�T���/���]�r�RU/���t��t	n	.͙��ۛ_~��~㜭��ٽ��ZqPl�������{ /j<��X�� �N@�M8�L3�	ǆ�
�]�s��I!p��դ/�R�v1��\��ꒄsC��;m�/����N��t\��|���]�x�������]\Y��������[{V�A�e�����%u��Y*-�%�!���ڪtMV��:S�݌�=�)��H��ϡ^a������	�?-Z�'N�k��dc�f�ZFHajj��}�S߸���}�؞?���T>�����h܊$P�v�������uwt�#�*��R�;�����j�WU��r��7vl}�`c�����6�l�FF�w�)�f��f:��8���q�L�PT̕���	�ė���(FQtt��D����_��7d��R,���O��XS|a.��*��R �/%b��ߠ�iG{�;�0T ����0�,Uy���|8ױ�~�!�X�Z�CJ~�]c�w�(��j�]��P��E!uL�b�A�ė|�������Kgv�G�ȶ�~���yw\������O~e�N:4��PT�5H--m�T��g�}N&/����2֠��:)i\�6�)�F@�(LKo5x	i+�4�Lt���+H?�N�<ϋq��|I����j�k+#���֝Mh��B^'ߥTp{�p �eAW
��$�H�.z��>��i9�jߋD^���*C�,���ܒ[e�XAI"�Rld������%�Q6}���� {;��(�g��8�����G7mjf�Jw#���F
+kC��U'%������4ŭ�3�1�q3��nu��^����{�0;���kh�/}�-�x�,D����U{��K���l�U��j��]�����?��}�˯ک���G�k3U�~#@�	��o{�G/���0pau���l���+��}u��0�+P��i%uMtDœM-����b]=����oKӋr��C��@�G��G�) �2֟E:�:�����5Ȓ�B��rr�$���cN���5,�/e�aai6h�@�5QA���W2��~5��"��(�1e�BD�HE$�EnZ�su~Y��l}�]�tF�E~X�3幋>8{Du(��N�ȟd"�ყn��� 4��L��6���F�!�W��y�&T�CZ�$&&J���EL�8�i5��y��ISSXo�#��N�~���;\r�vK��Mə/�F�L诋�;�X�Y������,�YvAݲ�Ŭ[z��f�t�ܳ���ʺ�.��))AL�����ll�k���W>K�l���y��_���/�}gw���t҆��ڃ����a�)�WG}/������)ZJj��LB~c�-���:����xP��7myE�V�����/Hp�]9c=�mV[�� J3g�Z�"�X(z��@� =��.O|��ΐW��h�H07��b�F�$�ʌ�
l�J/)��P˘��O�1��Tn;�*Y��3}^`inb�J��^{m�ҕR�T�>�X\#��$G��㜛�7�ǂ9��R�+B���2�ẘ��8��MR��uCK�"��b!�	0�ⱸ[| v���`4���Ex�t'��BM,%�ک#���ή>H��;67Y�:�+SG'�lvvݮ\>g��tZ��*/��dce��n&ȅ��0�yBq�U.��,���?'ˇ������*kИ�vX�gdȢ���Չ�V�q��SS�DȶĬ+R<33��$Fe��|���1�a���m��>���Y[Xҹ���`s�����f$�+67�dc�'ldX�?���z/�5<�{�{���ש��]�Ɓ�6�9�B�	����[�'��:2p���B�f|!G���B2��D�-�������}�����:�z& ���T�Sv�������g�����U;u��^� ����ǟ��k�kon��P#�.�{�K��_)�Z�X���ƕ)�PFc�"��$
r��4NX�YU�4��`_R�6�.�P�掔}��t�Ⱥ�{��r�dB.����r�/{���0D���~�R�E@
	�U��i.o���*�U��(h��{��<��m]�-�$a)��U��֬!`�mATǾzn\pq+���)��� *}ʤ��$͈���?���g7�(]W�v7?}b��[�;� ��,B������DW�	QmO�p`e���� ���3�~$ L����)�ױV�2��;��Y�-�^DĂAS/�G�Q[�RL���dB�!�P��Y[�eaIЎ�"�Rj��g��֎,�|����l.�ߑ���u��Zy[����?�R!����'�*��,N��\���:뽲�/V��`R�0M�����
k� O�
�_�#H�Sle!k����O�m���oO�x߷Bb2~zl�n~��f���$y$�W/���",:��+���S����/~�+�w��G��k��'?{�=�3h���ڔ����v��"�Wd�CO���D�j�Y�(������K@�����Rv�H�õ :�%�]�����Y,�F��Y�ǣ�j��w�d�8���8s�<v�������~ɾ��/�?��7��{�zz�u��&� %���#;��K���E�M��9�:��8�cAPQV���Dv9�ڄy�]W��C�l���-(��ڙ+��ڗ/x�ۆ��n�k�>{b?���6�Dᗐ�`����ʮ�����7�CK��R�))��D��@|����R1�h��0U��CK�+b�mi���P6�ђv<��DY񧰆,d���4nN0̟��i �� �ObKsB=J����Ye������Y
�w)	Y~VlJi�l��0�lBȞ�lkŲ�^�^�C��ݖu��]\X���{j��b�\��f�� ��J�6���e�틦g�mM0ujz�V��Ou�z�e���7m�ᴠ��N���$Lzj����z˲����<��ƀ�W%l��a�oq�dEQH��k�v����h�2�:1z��l��0�S�O"�{�.¾����fjg������ 9{����|>'�!�W
����]�9q���,���tvt�Ä.E*��zhR`�� ����G��@ I�D�<a���,F(Ap���`���zP�ϭ�Lt>'���¹2�D~��9����;��yh>��3��W)/����'���պ����D�e2���{>�O~��=z<j�Vj1]󓛂as�j�Ã��k��-�?���IU&�\���tu��U�&�OX��O�b�����MϪ�f��W��󐑡'� |�s�t�İj������Y�|����D�5�
�حe�@�&�� ��2j/B��Qg��U\b����y�∪�ˋ��8'�J3�����V��80�|_dڐ�4qHC�F!�XE�ں;��.��i����3:j�t��U��VcmR����n�Km[�u��]'[�Qm��5���v��)�M��~�Pc�*��X���7���isT�/e��_�Lcʾ��$�ORsRD�sV+�WߺdRT(^Y^T{�J�O��9$�nk qxQ�}SJ��'@�� �em����]+��1�P��iLu��ʨ zO�Lz%d����laa�S� :�KY�-k"�LFK˖��4R/������S������L�؇�����d+�Y?fܙЎ9���̊hB�.��0��s_@%/8�/5��?A�g/���`y	s�>����=s�0����36:4#�w����'���{�FGG-�]��!�T����3�K&���y�]\&?s[�S!�&+�`��[������A `3̆�M�9�bb�ڳP�"f��u=2�� z�מ��Vc���ڲ
R�����,|#,7K8�{���2��H9t��!����0�3�2u ,�Z8L���
�;��.��������Xj��������R�I��jwII�Z����׮�ͦ���A�Z���_��lm����ggΞ���v!�:k�o��������-����lW~��C�kI������>!�F	ަ�^c������N��J۝OG���]/!��g/\=e�u5����7�פDq�x򂄆��bAS��El��U�ʼ\�	_��nx�?V~�c�n-���#`��,:��Ю���xh�����P�/�.Ã��>��d�^�W��@;R��(�`fJ��`Ԇg�?ltd��?xl2F>H>���1N��L�<�(}����;2��0���<��UKs��)�S`�Qirl��gsm�F��û���ç�"�6��`ز/"|L@� ���$�ε��A��������,Ҧ|Q��������x���:T�� F���W���,�21-<�i6�{�*h��&A�e&��	� ���O06im�h(#��5+���̪���	���i#��+aF�������}�Ⱥ!PD`
Tṏ�L��	��z��Y�mL���iDI0�D�X�lg_�]�x�n���������ܸ���'�����M�ۭ���)!����l��s)�9}6%�mB�Vm�&��g�\!��B\$E�0��u�"�� I=���~�W���Q�W� B����ܔ%�rܵ��焪_�@�l|"]|ŋ1E������� H�F	�E��W���(�Gޭ��JמO+�	�	�l�1"v��<���~anY�b�"mmmᎯL5˿y(>�1�G,
��/.��q���2gj���fb���S)Ix���
�yف]�JLH([��;Һ�O��PH�"�f�!�ii�Z��j��$-]S.�8����Dv2��I�a�/#�K�(&�E�#�$gV���N=!�H��x�@`^����G� ����ERi�g�f�ߢ-��MHX���-���d_+��4G����{f��C�7�Ch�-� �l�]FGK�Y�D�����w�{h�}���[����K��̡a�x|7�3�rJ�v]�� ˹��5N'�X�u������G�N���O�,?���:Y���>�bu��=FFƄ�&'�������Ն][�!elE
<!ף��\\c���oS��\.���aˋ)g���lt|J>%�
6+��4���ݻ�@`Y���j*���N�P)4%��K�%�Ii�׈zVH�V��o���]4�P���u>��A��ox��0ь�����A����s;;�V��MS|E�]��.�ie�"�RE��d
�)Gs_�y[�ݕ����9�p-�5X>y+�����k5.f�%��>�Yy���� �C����tyy��훿�{��s��V���w5ەW.XkG�[�ήV;}��.������A���(X�/⢕��G��ԋ�)��jVO��Ղ�\H�fqa�J���I���ߛ�,d��6��Qj����p/��BِEC�ur�x�}U^!��$�<����]��T�8T`O��X$e�P�R��a>'��̕�,�I]ס��Gx&\��{���ɂ��WEyR�T����<�sY�aK�WX�|��|���J+S>1��N��v�)������Ԫ�����Ox$a���x
�Ndt3�U?���2���x�|�54Wj�k�c���O{X�|�T��kc)��n�����'�t�-hF��&��eV��N�B�;�cA��C�1q���(�],���xŃ8���*|q-D~�������(C/�C�$��
�h���cτ���C	�@�yXA#H��@��`�_ FŹ%���	�*�����ϸ����t�k=M�4n�'�;��5����Y]���f�7�qD�L����͚�뭚��5`�|r�W�"%΀z�����K��l&��ߘc)+��v.TX�:V^��@L$��bT���k��o��!�cO�]����q�K\��m����BK{�g�PZ�6��H���[�<�B�e��֎�;�BIȣ\ߕ�UXUu���Ё~�t�x��������'�汲hb�P���(�4�F���Y�}��gl��=��ZD<�AMU�ϐ,L>�oD0P&S��6h�7lvj���*�X�h���ɰLLY�>M� z�~'IAʺ�j��a=Y��4g�C
�i��t�56�� R#���������M��K���Xa�	Ԅ5G�2<��g�A%PQc�R<��~0!w����w!�n݀�>���¦�◜L���p!Ò���bO�~0��ȴK0�sm� �8�Ǽ8y����ɨ����u_sC�w�K�C򙋣|��$'w��L�M�=���j�򣶙���0��b�d"-�,Bn�-ήؓ��4���m� 8�XV�Ɓ�G
N� ��	� ,.��$�G`�k�q�R
�K��uf�Y*|0�E:�d]r�+.�M���i�4�ֵ��ž��߲o����k_}�:e�W��=��LT�?��w���ڹ�}b�a1沵t7۷~�%;}�_>��k���/���K�b��2F���r�~�G_�&	���q��^q�C1餘'0��9-Kw�}�/k�SP�D�Io����OȒ�3��]ф @��KYу]xlxx�r	��)�rO����
��YeM��,mm-Mv��#��y��;����FzU�z�[��.�JV�B�<W���Se�M�S��v�YS]��~�������ڊP� �{��<E$w����LJ�h6����P��L� �o�%�����\kE�7��L9�`&b�H�씌�K� ��h�k>r�-1������7����#l�t����4T�	hU\Vd���έT���	杙������Qt>����k�ˮ1��,��e9i[T�-��b���{YIV����q(�MY/6^#E���g�]���������-�m��Զ�Ni�fi�Fi���A����}�"��$|����ALɢV����k�aF44n��z_��o�f��������ٮ`��-��`�=*��w��Ξ;e�5�V[��Y62@JJ���+W����V�W��<��.�]{�mI1�V�S?{�;����w��ׯZSC�MON˪��W�-	�[�_�G��|~�Rh555�w�ݾ�����?�������ׯ��OZcS��MN�#��h�jt뷑gc6�tT�&�1.%�o���������Ձx����g�Lw(%,h��GDO�ꖦ:���Ƣ��J�7*�H$���)���._9c����nŨ�I��C	�+��vM��ή�ٓ��mjf�gu�u�y��|C��LV�%`$�	���G�o��5�(U�,�/���(@p��5�i�����Y^��[�y���Q� �h���;[�O���|�Z�-�0�g�%Ô�D�(�C��Y��70,���o��L*�C=�y��A��yg3����M���&�h��g-Vq^�]���`�r�s�8��ٚD�.[]��]#M_#%Po�Ui��Z}^�������\��ϲ���梬\�mot	r�YE�Y}׫����`ĤHrtVH�H A��S���r�3&�	ӳ�(#�~���_�zOv��~����_�is��Xo�ݭ���f'�۬�6)zDc z����4{xxth�nK�N8����t2� ?x��߶��z1b�4������>\��n�ݰ��}52��ki}d��gZ��YY��~���eW����
�(k}]�����g��l͖�s>���C��U>�h�a�MUv�b�u��x��DU�N�ٗ������Vi���=M��F��η�m�wA!�O�շ��7��O[K[�`q�sϝ�Dl֘��z1��pE ꘛZ�]7��/���-����/ثR:'����'4�>����y�,,'���$�7��nk|H  �<��0�DJj�s')�
$�y�Gb
?�0)!�ꚴϥr}������� ݉�r'LI�3A�?�H�t�j����%����ɟ�^]�TL�Z%��S݉����&I9�8�;�E+;mU�I��ʒXe��N��sʒ���>1w���&�lKK�65Qa�1����1����X���Fmb<f3SI	_�,F����%b���{�,�'�wB����>Y���o�3�@��:�Qj� %�`@^��m��������$������81 ���������ɫ�"Y���2���e'Nv�me����v��R{��h˦��Āܗ$B�(f>���)��9&;��FB���@-����݂0}�Jɒ����qA�1��;����(��z����snE��Ro�^�ll�����W�B�	"��k�l���ŘM����h���c�O�跾�~߷�^�Ѡ���E7[ks�u����ؠ��+��R��ljt^�r�'տ�;_��:�T�J�*�86e�sR"5�)� ��̧����)������˓�#6;�h�j�I	��K��U���<�**����j����H6��|��,�E��{ҚL�xtVB澼���W��@��Kdߔ]H�A���	��Q#y���EZۨ �떆�+6�v�A'���GbUh5�2$�$�-����
L��Vz8�P��+�)|�
��uߝ-�q� ��jF��Ŝ����gU�S��ye^�kY� M�H��[m�����ݷL�e2{H9��B/���y��Ӧ�l�f������{%�:���qC�^16%�:e�� u�`�GEd���� ����o_�����}U���ىS'�Jд��͚e��>nH�M�.���EY���5[Y�v���X�!����͔	F	r��ѐmi�XY�ڒ��.�㇃6��wŀ��Y�\c>|0j[��ڸ<i�Uzά��,���oJYOO��o�:��?���{�jj��d��,y
ܲ�x��ږ64����Ip3��5�2�9{�tL~︔�SO�}�������a{p�}��#{�و>l�n<�[<�������v�����}OR�>{���"�;D�6
664�֪�����.�R%zi��i��P%�O&�٣q_ z�b����+Rz�&��n}��n|<(�4d�~�@(�D}���%�V�VI���2�������/��9!������
R��)��*2rd����Y#B���#�Mm�K���d�=#k��̫07����`$�ʗc���,���{�b2����
A�Ki ��/�2�[��%ō��t���ڮ|iK>%�cݽy��e����n�Đ���|�i�8�ag�l[�~��嬷7��6��gEZ����{�3�am�K�xC�w�P����Ufm�Pe������Ԝ���A���%K�)g�?�9YY�w��Y�듥5&���ٮ/C![��sTȝ�_�6���1;P�}MN����c666��K6�k�%���ٱ��5�����DH))A#8�&bG����YS�|��o�&��Q�))3|k�%IЛE��q_^���ԊO�T�A��dW��Ҝ��ִ��e(i�7u��r��L�0!O�̩����5)�a1���1A�9[[[���� <���)����Q}?jsӲ �:oJ�~^t���/�S��=�-�x��N�W��ߴѱE�66��1	!��[�+316g�|���&仪�/�zA0��}n�*�w�=�5	�,8�:���`��؄h)����#c��b��}>��A��TnE�����uG�!�R��F%.�����e!����p1�Z#8LL�ؐ��~��`>�+��v!�˱C�+k*|cn/�#�$�	�D��d�gN�Yp���|����n�r	�:�[|�R�Y��x�������^Y��E��fW���memI+�&��0���?����?����U�t�����u{��v�L�`Ҭ=}�̊վx��l�AD������Pl����؄��d�	1�N�/;8(���6/��LUK�f�s��a�TW%wl�D���o��l36֤��ؐ|���k��07���JAB-g\maW���4?��Y�D������	D�G3�)w�%�bD��'e�I�aA"a�q1�` �;�J�,����������&	��TE�<!���Ir��9�p7Մ�W��k�ik��$%"�˜Uq	Q�m�V�wkE4"'��P����)r+�R��K�[���͂��EB4����Z4��/�J��XgW���V�6ihK[I\6K}�l�h�n;�����殍O�Rn��^됿]��w:�?��Ħ�'%L�<)T�K���ǫ���q���+����,6e.��
iD'=R��!r�򹜔/y��sIЎ��v���О���t�K�Tׂg��������������'�ł��"����L#�B���!T&�}%��,)f�F_pM�[���[luf��_8c�N�{�R�a�OTF�K����_�l�b���zi捄���W���Qb�j;s~�Z[�՞P���g��xDV���W#�,�0-&�.�*&��� �:����Y�@	�(�b0|�Z����ZK�7Ś���'��x.��S,��."��j�w�}>��e.^k�)0��r��e"��B��e�i�C�ӓ�-F_�X���j�������4l�0;�ոF%0����&��w)��^䉢����ߏ��2G8�
6/�bWj��N/H)���v�χD��O	��?��y%S �=)�����	�4X�\#+��!�.����fi��D|�ڏaJԯ
�ͺ�:KU�l]y5K���ۈ�;�4o�m�ielX�0 5$�8)KF�f���,�R�a|q\�P�Ρ)SQ�5���Ke����J�44�t�f�;�r�):2�㹤�dM�-�	
�E@�mh�v� �Et$���0v�g�f�l�"�B0s^��p"6XGB��Z�&Eh�w�-����=���l[���������lϪ2ID� Z��>�g�����$!\4,U���DD�2���F�����5iiv�l��=�!Y�XJ��T�LB��9)��c����oE�"dbA- ��l��܉(fjlk��Ҡ��E%LV���<���E>GveR��h+�H��6::'� ��L�݋i�X��.��4'rU�^_۳��|�e	�=�|8fCϦ=p��%&����F�41ao�L骄�W�R�Xiw��1	O��
��9��A!�y\����bhBtf�����ɛ��w�a���B�k��Têb:�� ��B='��R�M[�����3W!w�EA��ڍUF��75��dQ=�D��r�����	Y��8���S=.d#�j�e4�=ƝyO 5�b(�*	q"�dPX\�;�;Q���i�������}b�'��A���@�
갗T"Z!���Kc4
6�w}���XM]�����#��
�0_�$ T��iK�40+�R�䐖'[�
��	р$˖J8��iI�{M��)�P�=)Ky9�k�&�6� |>�n��[���A��k��mM�+l[���Ҷ��>�L�c�\K��� ���>��d-��9�0�F���hР/�M��aH�aP^h\|��3H� �.�S��m�K+���df��T��<�gg/���^�^z�5��[	y����J��'hV*�^l�1���?��/\�K�O�Y�3g����օUu%G����@˟�R�R�0���⩢
�1
ㆵ$EM4�d1��HT���lmͩ�;���!D[�����,u��ט*��K�x�	����}r�9���Qb�� gi�� -U��FU�
����!ᠳ�E��ǷF|Y���9�=���-�O����Ec�~/�^L� l�nEBʜ<�ꪴe��!e�b��`gQ	]2��YMuڣ�<;������ڭT���M]+y�{Z[�7�R�.@��놖Gb�Ȳ^h*AP��Met>K4H��O�+����W����	gcZK}�9��}i>���QJ�����<�*�"�D��Qɭ�ze�qF��U��s���鈴gZ������X��tn��FwR�w�/&+Y�Y��`@��0����"��To�������@�IR]\���bSS+TB�x�����*{�K������&k�s�;����ɺ�[�ԹN�x���#?o��.\��ﲓ������:�Z�y	]'�V����#��\`,��x�#C�V>��m�|IY�P{?Xlg6i�B��<]�P.�-���*���(���(4?�@���"sr.��q=�\��fo}񪝿xZ(B���p������$���x�XB!v��D@X^��d_�lx�"%׃�f�F���Y�q�{���ʑX�� 5�j����}�cI�f���@�u���	n������J@մ`ơ&
Emq�GhE�+��S��\E�T�G8���X\p�<^�~C�^T��W���AL*�+�hb&Ү\��Q�*�`�Je`(��G�ԎP��f�}�K/[{k�C+��z�m#�Q�ېVc&�>Խ�]Rl* G3Q��N%��㘛N2��9yF�M�4�ۨ�;,�o_"`�{K?px5��Jˈ���j���0��n�#���@C������TӪ��q�g��I���*+�/I���Qb��,xQ�j3����k'��|��S������v�<�nk���&��2�ER~$S_����E�͊���L/@�n)A^R����Ȓ3����/�^X2��	�~$���B&��� ,��H�`�HPF���ܹӖ���{���H�M�I�"��%k�+4�m�0lm��ZN�r��������$�c���$[��V��ɒIaa��gjA��ojZ�9�Y� �$�~'����&�W�2�R�Ȳ'΀b�Wı ��R���{�/2�$괬+r�W*]U���DP�}��Jp�����Bє�q�˸I��+#Г�'ՇK�I� X�y�롞����ap��;�v��K!������o��`���4��c�)�{�T,���k����Z 5�bg�����X]��{1+`7��38�AC�Ҷ"ע�=�J���Rh��G�G��x)f�������x���1�@FUu�K��97�Ҥ	���J�b��ZG���K�J[JT��h���!0��P0�)�$-@�ā �������4n��R��	�Y����&Jw�=V��DC^���
���qD)�]�.��� �I�s��V��@~���xr�7��R�u_��kټ�ꚗ�#�
ߌl�F�x+��j،�C��,Vr �E|)(Iy�2�QV\�bAsV��^��`�N����̑��gz9�����H�غ\�-��*���HProS
G툆���b-Y$��{Q	B�\ZcS�]��i��vXGg�5ȍ����m)�r�ge=uF���q����҆����ciZ9�;&a���ض�%�X0��3�p	�9���pD���T��F5�qr�X<>6e++k���JH�	�2�����e�;�����WAb2���²���zEl����rYf�UsF� �Qe����g���P�����Q>>)A bSV��|��lx� "I��3�~�/���+�/fLH�Uױ8UH��I��կ�L�9h>� 4@-
���!�)���ޡmI��x?����|:vv-���,�8����u���WO�ɓ�VS�ֹ������N�@<`�z8����Ɣ��a�P�T�*�����t;�#%'Xq�b�PR]����x/�@��8��M�Z�\QRn���ȷ���n�/��S���S���d�M�u�~,�%ۦL�o���%�vR���^���^R�>��u�~Y����&e�em�B���#����Aq|E�vC}�]�2`��q^0�ק?��T���`���c�����Q<��lD]&gM��ut4��-�L	s�dO�-
���1)W�9&X�p��\�cʽ&���% ���4[���*d|h�왵w%�ʕ>Z�|.	3p���oה���P��8�)\�Y��Ŭ0���AXx&��(7Ed&�O�������b��f�}���8ʵ.�B�B�^���+�� t�h�bЦ�Z�?F�8~�\0yO�ą(���S��U/�Y~U��9C�2��u��E�5���ۀts�[�V�5��u�n�'�>�\��:i}�mv�b��x��]}�]|��kT���֝�#~���:|���ZRYZX���E���3ei�����/!pX����\���وT744ڵk�+���$���0��޸g7u�u�����J9��L����L�%.+�C����)ʄr'El��M����ڰƶzY��mH�
��0���g�#ܜё�6��/)Q�_��jnkP�����̪�$u�`��	KHձH[[�;R���I�J@��d���*���O��؀����4Ȗ�L�8�m���������kx���3(��IL U�'�v\�=,��θ��ߡ�� :hS�P	��ܲ=���7�~p�=��Cc>'25� A�`HC<�)�,;<ˢ±�q{����;Ũ-j�,ߧ�_�E�M��B���)faB���@��A�T�d2m�TJB�i-2���Q����A�S}.�ǯA��0bKs�uw��*���f��$:���X����r�e܁�����f1T�\A(��n=��.�:&H��9!	���e:�*?7����J�8���<��¶����-/,����MO�:�y�L�h�PΠjbf��hPR��ߕ������yU��p��|�t�
7cŀ��OG��O��²�Fh�4�����B1Eea��'��ؠq��.�����!��Ԭ����t�X��>ߢw�񐞴��k����A
�.�QK)T��mɈ0��TLH ��r�������.d�g���$�D�l�7<!hc���;s#�{;� &
E� �d �4���E@;:M�'��޳�FT���w��&�a���|'@�� �`pI�r����fc���{��˟�o�}v����i ��;�RX���a{�ݏ�W��M>��ͱ�h����u�k���3�p)�(��b�����j1L�0%K�-#SX�B��̘� e�o���ne��q���@?��� �K�j�L0�T���n�tM`�p��蟻��jc���r&���8H�Om�/�Nʮ�D(,��=</: �<��?S�8L�iy�C�	 0���Q�X)���%��d�p�"ʤm
ip�(\+�����Ј�۰{|!4 z?}��>���
�����J|�l��39Jo��r�y���}�)���g�@��>ާ�Wz��g�Z&�����%���ɑ9	V�y��#0EԼ��"4[�6Яw���!=��=|<��ā�($*
����X&V���-(�I@�}Y%�;���������*x��!Tvyw�`�%���J�P���&�2>�����H�/t������2�:�0�"B��6�d�n\�̲�u�����\b9�l�S&G�<)�Ѐ<>&A��&F�H��[O�?��X�J��b9�u�L^Z[��[j,��K3�4/}�i���|�-{���2ƙN���@���*�3��Q3z�e
��,�0!����a��0�3�_��խ�9��s�
J �\�����>�ͽ%�Յ������g�źO��N���`!u�f����k�i���F�0#QAc]�\,��=��ӓϙ'u�H�)Y�_��������=z�ܶ�L+fn+?Ee���{�aqY�X*ꁫ�����Gc��3�����3� ��s)?�b_�lvC�FFAk��f�8���P4��`��r޲��Ra�`w�6
Y��e)R[ ��a��u��d�jUL8�9"$�/m���`��e˯d}��>�{w�%���(���B3����y6��C�hc���ʓLF�&Q��	>����WH?����ơ��,�׿��s��A�`�f�@����h��Mi�]?gvf����u�@����mo#�L30�0N8E�(9��{*��*�S���7�h!��(jMm�����Va�i�OV����hB���ǆ��?h��B̀"@0��>�����Ƌ(����wj,AȨV3����ρ���EX �1�
>�� a��E��q깏���}[O�(i\r��]ߤ�a�(=^`7��M1�|�<�]��6t�`~�,�����h(�j��mY-5����v�7ˈx_,�^-��;��J���@{��ڌ�o�7i)h�3��/�.�b�"���e2@sD��]���ʢ-/΋W��/̣Q�!;tm�;0� �a�����Ǣ�K8ЁZ����-�/K�'''��>�?�?����߳�>�=6�� ������u,��D���8�@��¢�d�?���?qQ~{��|�� ���R����>��P���y�h"�O'h�����<��R�bq���1�g��7�Fړn��� ���N"K�E	T�6�2���^?�͜ �ک>�2�֗��+�A�o�%ttr��:��R��H�3��&��`W��������!����H0N8��u�ň\�!����7����t�p�[ &l]�����p�PZ��� �0Υ1zJQ��� �w��-�󟐟�ڭd����~��R>YI�����'2�WY!�얕��6(	��JqKBx�1=c�.X&�]	T��)�����LR�h�/eD+գx�#�OJU��^[PP,W��� ޲Sц[�I;����k2<�٣��/�p���E��)%6�������؆zY^7��C��I�y��ei�I���e���6:6���� E9��^ע��˴�Pt][��9.f�IzN�"a�$���G1�0�^�L�\� 9r�33>G��|��3�s�_�Jrmi9�g���mYq+���# ��6��o��t8X'k.af*{wE4�Q�����3����ݻ>��ǖ�W0��-<��+ƽ����z��3٪���
:&������ϧ�>��w�=/���N���4H�������t8t4�=eh�Gm9G�b�F�{��s�]FH�V�RL�II)������pO��"��Ϡ��ú��̅�'}`�2pᑠ�C!��b�قf�	:����K �����ó=��͓(��=�4R<	b��j���VW%�s^O�=�00��d��uy�ł|<��\��<H�tm"j�9���YρOeZE�55>�F����|UR���"I8��QA`s)i�x4n���:����Ģ�<����5��}4���h��� �Dg8��"tD�� \�Q�sbq���i-�+&%�Ņ'"�]4�qp�Cd_\���#"�Դ�I�QK�(A]��8o�uվ��W�OX�bߪ|�$���pfV����^��\��c��b��si�Dh��N����s��u$T|��p�S�I���N
���e��0f:���0��g�u�﹟7H�������/_���x�+��5e�H��*�$lL�����ߖ����p4"��[+�Ot<�'�8j��*>uz�`������u�`���E���P�E<���#�x�DL.��{�+���0<C� b�Q��!�O�˒��U[��Z�X\��-ؼ�y��s�b����t.-�laqŲ�5��UY�%�^��%���_�x�u��'넘�yWs6�t�&��[n5�2�%�9��8*���#�(4r��|C���-#"�2к'�#�'���a�(I�������u�<]��ȖCl�4��#k�3�D3�H{�<U��W^�����;?����ٷ������y�!bb=��1��A�@ԙ_�y/`�O������\��
� m��G�ޣ>����A'}�{�r���Q�r��;ц{X�e��GGy��p[n�k���K�d:�f۞^�֛/�׿�}�;_�o�M;��W8�M��̸4��-L-��ļ͎�����^0��͉��2z����N�T�h�����h����-XS	ő ��0�Nf��P�W��㸞�)�@/O�Kcʄ��-Y�	u#y�L�ʘ[P��{��X�NN�@¶"�$e�c��D�Q�'��3W�1�H:��;�$��/-�ɺ����}i5���H)$�9���؞����MOH�)\�c��nnbkPuL�y��\_���X���/7�h;���s]b`05f�zgD�G�8� &�Ԥ��[}� �ׄ��Z��X ܊&z��#���}Ѿ�ŷ����R�5��ci=[m� �.�I_��!|��6�C4��ʃv��g�a�{����	���p�C��MP.��h���@��=�p�_���-��AQ?�?8��i'��&��0D��Bl���ݳg�%8��,�إ�$p��ŋ�R,L<���_�]c|��	{̱�(
�]uf�mR�ܚ1��o���*��ߎ\��η���D�)^C?��F�ƃ���ƪ��J%)&�Q�,�a�����w�� �R_�BJ��4���R�L�(�e�H~���n���q`�����!P��L�ǉcr�ʾ�a�j���zx,,��x�h���d��Ҟ���2A��ks���3p�A�a|��{F�`\�����fjǱV�3~�. �
ͦÙG���2�5	wL	6x)6��8d)�\��ܓ~��Tq9�g.\�+W�Y���� "��f��6/M=16��J�t������_? ��F1�ڌ4`oJ��N �I�6r��ڣs� �[�����#��&�)�㧇pc.Ջ����Rˎ���x6��5X`,m�E���!��gD�8�IY�-��?�m?�������Xgw�}�[_�g����|�?��胁��
��-�� hN[��й���7��cu�����Q_����}�g;��O��l��}�m�z���.�^ԡ�~�����͂P���1@�zEF�¯!��7��K���������PK����Lx�����G���,\��he�ˤ)N+jDI�X,P#:T]S-L^���V���HJ�:�����>���)kl��À)$�rN�Y̳���>BƆ��\#SW�Ko�V�3� ��Ak��0�k)z/�} K B���|�S��KȞp��g�����d1"e񔵶5���C
|L�wG��g�	b�z[��,� x�sM=a%�f �s܁�$�X� � %��O�x�C��=T;]`h�ԇ.~�S��H�����-�T��]-Q��T��Lm����<n�M�`GB�sxωN@|]�ڸ�StWV���{��ڍ[�m[Я���Z���Ø�̍�Sq	Q�O��П�u��儵�PS{g�WP�e�RHG��1<�}��I �nw�u�%�w�Ú��u��"��O��E�]a���f�<h��D�=�Bi�pG�P����r'�z{�@�P�f�Vl�鴍�
�,{���X����?񪬊 a64ց��2���e=m^���Z�XځN}�'H�DKvݖ�ٖV��®��nK��m#��10rP	mJ��)��=���0ky�;D'6е���C	I� {!L���>4�J���	��A�"a|��z�š�E$h܍��hu��wH�N�wX�2!�0�m{{�6� 2�7�HG�|�y��3�C�a� �Բ,ȿd�(�hp��Nr�x\Wp������Eh����˳D�{\�p�*��uĔ��hJ	ڑ鳺R�����x���И��7�+4���T��������YGG���Ǚ��}N�10��]/+m"R2���^g��tXL.S3�4�� l�~t �
+���`�/���)Uː[�M�C؈FR����J�AUY?����-���B`@GP��"��S�,�*����Ue�B?e^�>���g��@Knu4�q}�5��XCK�ާuYi�M�K.W��jH��+AR/5寿{�~��H�S�vW&:.����W&Sΰ���!D��ֈH�M����>8�*-W.����W��LF:ù�i0D�d��K�Z[3�a�6�D�\��gXb`V�1rR@P����Ɉ�b��/�.M�@�C��%~#�����s�\�Qy�����	{�xʞ<����(�髫��`)��{<��q;���P�荥Yj?��eG����;8?I�ޢ���=�e���G��~����������}z���͓�Ki�~���m=�ND��%��U?�nXs�`m���ܲs�q{rP���������$H��W�Z_z�]��o����^b!�?�%��DA)�d�=�h/�~����2w�'ƀ'����g��s+9+�o���b�YdJ=�FI
�?�f�j �ik� K(c��B㖖��ZB��0���tB����(ypr�%L�m�2�Hu�MFw�v���h)e�mQ�P�p��r�������?)�B�UDd�����8M��Shԋl���%��Έr�5H�xxp���4�{�li���_� �X��+�\���N}�f]�VV&��=�N	�ft��f�c㶲4�{���������M��!��skv��C�������w�?��>�𾭬���������Fgl���?W>|�m�˛~d��:�3�K9`��m􁇪�<����G;%��n߾o�?�g�Ϟ�������̼[��{��X2V_�L��	i`�	j0�k���9�V�$#�hR�B�Aۣ���#�������K�����J�C�'��� ���Ɣ�p��^}����M£gHh��+�HPD[�,$�"��=�������kcS�t�Q	���W�u�q-�L$�pRMU��=I鳵�Fv�v6���E��/b�����E�2LѸ�T���!�(��m&
�)d�a��u_�-��sC	�4�|����b��:x(��2�-����Yeʄk�d~a'�^0��C;�\l�]�,��t�׾��]��)-��F$�+b��H���H�Ξ뵯|�Mk��V7�('~&�롥H^|^&� ����K���E�����*��6��6WE��Gt�H��D�"X0���� ������S���&myy�Wv`��D:ݏ�=�1�����v�Ac�7>�"��=�u��|�4.X.m|�U0�g��W��A	��\Q�q�H{�k�di�6���Z�'a���XM|�*�d��(2��i��bꅵ��ՠJ�r��t�b�aHJ�y�\c!�Z,�������i_��+v�k�XS[�؋����|�{镫�)�P��'ӽ_��`��[���QckX�}�Rr��8@N��<ؾ���E�=�x@VƇ��Ϋ�Pz�9�=�^�O�}�h�����x��V4�,NP"(l��Pg1i��R!�QQ�JA���¢,�FChh�Y0�^+_?����)��Y��x��X�3U��c\�cC[��ܖf�,�h���::�;���}��o���sd��g��{�t�}�koؗ���׶�*�Pp˗�`�h���s2��@�X�Jݐ�Z��z6ڟ
�,�$L�F�q+��G�x0Ў����6b^Y�"�(lI���RFA��O,>i��1t/~�>��GMt��5���xv`l]��5��̭�]����X��EO�,E� ]-MϪ
ɫ�ϼ�o`%��`q�O�/	]}��~��O�Jfw�D�+Q��TH ��h?ʃ�t�Mh,B��ȯE9F|�^uU��9��W޶���7�?�-�܌p���ZyE��	r�J��ׇ�8/���dA�������&�_!��W���3��b�;��=��=�xeR�aXIP�bv/��d|	���OJ�CEr��ɒI�h��d-N��N�&���ܤ�X�����f���b+��-�"���.�19�\K)C0L�����Z͵��HC�V}��!��E�E������w��w���c��~�����~����׿�����>	Yi{YJ�Āxp�ˠ��|�3%D0YC��@x2=D�#Pbmm��M�����8K��2�H�I�00_TZrh���/g)=O��S_a���#|^�-��y��3�^>^�=7�b2�K�}/�;-����Pu�GҠ?�D�4^$E'*� j�tk*C������3Bν��T�R�������ڭf¢h��X�5wՊ)��GiNRV��}�Om���ʿ�J�m�T��7�U騖����j���J��d ��*tt�BIR�'(1(����x���a+�'$P���$���Q�=DD˭�����ڳ��R���b�+hbXk�J�)�gcSƨ&��o�ϳ���낊"(5�����^7�]L���1V2��OI������bL�%��< ���@IJӢ�Wc娅��;���t��ߤ��$���b���ݥT���ɴZ{ۀ��wEE��s�\<>�1���K@d䩈LB�n.��Yʮ˩t�!P�0%J�}7���;���K9��xX:�EIc��u��R-�<���[���On��uǓ���ȧG�I`,)hH^(�����X����0�T�$]�����Q�UW84������� U�+���F���E����zߣ�X��H�,��c�
   �IDAT�{����Q6A�e�}@��nk� 2��І�H1k&���2�[�v�a(/���'˅��',ŢV
I��+� k�[6�l�>��8�X�pMƿ ������U�R���D�V.*!�M�;�b��u��S ��yvDV��gV� �������e��Gx���Hဦ*eV�H\V+�N�T</'��vJ�^�<�B���];X������UVWxU���(Τܰ��V��j����$Y��A��`l*G���VQ1��(��BSL��8P��dP�͆��@"T:B�)�Ԧ��]T����\�GW��GJٺ���p'��2��B(�"�Ѻ��2!�>������j���NA��A���tl�=^�XݐN��7���@���!](L��]�m������<�:r��$���})���	�}�7W�8��G�0��\w��G9�/]�]���q���f��f�嫇�].�eۦF�`��s	���9{z�>����H�ED�J�(�
1N�V�*�mYXK�t6�L`?�o����>'Ǘlll��	I�@0����rB�9�"�~�Ƙ�kQn(d���sO�'���WJ�SFh�A�c�Q ($�-�s@|6}�C��qYy�� �K2�=�y��ޒ4��6�� ���ʔp)��	 2H(X�E'c1v�'T/mV,���m�IK��"��TAQØT#�fW�OX^�p��0�u�!h�@��!#@b��Ä�:l���0p��H&F��ɣQ��'�RB�ף����:I�nl~vޖ�rb2�)0����rl)��ٸ�X�8�_���KK+�&)&�8�]͎��Y�<�F B[93soC"�>�����s�bq��}�_߹ x[G�K�q^Gߋ~�]<�
�>U��ND+A�~�ڌU���Y�[]W#똲Bn��{���!������_49^m�.����#��_�¦'�}�<�S�U7E�U������*c^t�!S�ߕ��E�R�/ "HD��M�|lx�6s�ð튛�b6�����z�Y�U.����`���D$,1���炮��h�������b/�x�N�YKc�?����N�%#�(F�bS��$�Y�0*"��h��ܼ,L'CC���o*-#��`n��Y�2�ns�6?�lˋ���򚴈��:���E���][Z���%d�bL=�+&:�op�v�JCX+�\��YH� :`���[�lj|A�:��09�0��G�ٵ��Y�}����*���}��ήv�d����X��7/�	�#Ce�, A�!�E�?Xh���@a���X/�v!�}�'\N����N��g��u�Ho��{�r(5���ob8� eꪥ��(K���ht���j�?4
��z�Z�^�X+8���΍g��7M^b�̢?L�,�c�PDtݓpoH	�B慧0��l��Q����UɤRV-!����%,��	VH�I�:�;NTȟ*_�{B""�����M��1m**޳�j	@m�S��J��D6������	YT�R���60�~��i{����~A�+Ћuv$[�;���o�=�b�c�dj��I��	3_�Ծ��I;}���[�΂Q;l�m��y7�L�b��]��e���_ÿs��r?G���%%d@��" Q V�2�6�D�c`]Q�l��NIc2._��J04��M��#���G��&a�Ղ�D�$�U�4����8_:#��a�A���rG�Ǌ5]�.ڍ�>���=�l�_�(�\��}q�E<�	�Ǐ}�+�I�����ʩ��e��v��Ȍ�X� y>	����H��0H(���>_T�{����b�B`h�F�����P����@$���X��MA��������$(�V�eZ���D�h-_��I��������lqyQ��B�Q�(�^�B�����C��8OL�ql�O
��g?�س{3��֘ڒ��li�`s�y���Ia��У9���w�'��}��N�FY��꤄�B�>Q~� �cԅ�q%W�6|_��)GY��&O�2�U�);y��u�ux>/�:c�݄,Z*����U�2-I��6�OT�
�	�rm�l�\�HW{�;�|�����b�E��'��t���x�9�#M��b�鸈��E/1��I���ܝ�=�YꕛX�B���t=i�C|ٙ}��f��t{w������A:A��b����C�	�"a�ajvAq�#���gliC�hZ����oۣ�Omv~�UՂ��uÆ[7�<���EZuC� yI�
�o[ss�55W�`�ז%([��=�ʵ.9}0��|��g�����Q6E�R�?w6�1p�ڡ�T,L�hA�_�	BsĄjP��Ap`V�̯���� q�c(M���P*�����trl�n�Z/-���
�b�PN|�T�;SK�[�� ��6?�`��'}א���v�����ʎ�����}*ڬ뱲�bj�O@D�`=��`��wU{ر�R
������:�r'��o��w��_߰��1~6�k'&���)�LbblR�}*>|n��9)�%zG(�����ew׬�L�����RUج�����_]���>	?�
4Ba���V��)��R���qZ�=h�]��e���D���̮�8��Fz��!4�v�����a���[��XR ��n�O���Y�0�����A}�ΐ�"RB��[f]�>(z�ϖ�岔���T/�Pa���G�޶_��|2)m��\���yi��͟ߣC3������G�4��8��MY��7���5�tY}�Yل���e���A��p��3 K,<��2`(ݼ)%�Q`�BZB�Ԣ�6�%,����@�n��L}g*15�����w�y��l�-�<�o��G�] t8�DP��`�~!��n����{�S���)�ߑ~1�#�y�!�ѡ	�OCbJ6�ԗ��Z\6�k��ԣr1"w^]���-�o�"�W�ȳE�����}��MAv�+CiЦ�Hi�>�/������n���2��ƗO��m�'�l����V��记�θ���Z{{���TZkk�O0��}s[��ⶰ�d7�?���F���N����5��٩'�}��r_�'�8�=�P]�
JI�T��!=z�@0  Y?\"Q�->t'�}�ג��ɓQ}&~��q��'�>�3�~��9s�������c� X RF�����COo�����r���٤�3�:Q냽ti��	.zV����9�bj�4I�e%m:�4ƾ凖�MfU�Q.��i�5]���9���5�О[28�8��eQeww��7�b�M��L����mm�@�X��Ǔv�ΐ4ͦ�l	�n��o1���#Aڜ�E>�G���0,�y�����=6e�k�M[Y-X���ѓ2����������T�X���b�=+Fi���a�Hᯠ�9�p�v���K�.8��<��A �5��t�	�ཱྀ�|��Y�qY�u�ڬ�b���
Q��*���6�� LN�)v��j����ޔ��x�>���0�!�u�%)�Q>�;��}1���D�'��G����!��/J(���\b�.��}��5g,͎6B'��M���YRnS�p<s^�O�����{d^�-���y:�w�}h}�V�g�������zcI*�"U�|��E��&�s��tr������_��
feɄ¾����Y�d`.�I��=��1!��h��g����rN_���w��!{ce~Y���a���Pf-+��_j��4N���ab��FΫ)	N����<%��.�]-���ٯ���ý>��걃�	a�:�j�KM�[m��hS[;��~i�^i�f����G��~��[�4N�wN*|@J�Iϗ0�N�8��lvs��@>��ڈSca�/�M�3�䩙_���*)kY)!shA�K�n��KӋ���(G�
�< ���������� a���`�?���v8R�{~�����)\rt���ӏ����HęËYSKJ}�D�B�xJ�2���U4	qT 
�S[⁜[���e{�`؞�Lȏ^��ݲ"��Lj3��+��5��4u�?V]U _���=3��/[жT�B|��V��5�����/��?��Ac������ZiM
-X
�5L�a�=s�����Ҟ;瞹�����k���Z�鐊�nv8?}�����:?uv&{�W�棿�SwĽ���b ���!�n�֖�&���9)��sX&��K.2�ק��¾��3�Ϧ.M"�Q�J!�6(�B��[X\�=�ײ����9���k�ݪX���U�ڻi+� VI�忼����_��;� ۶{�R'�LK����i��}����r�cc�bO���y<�8�@�6p��#�� U��DZ;; �����Lͱ��KFʮ�RxyC~I�I�Ҵ+�}gA��By�B��#�!I�2r�ɹ��;Jyn_�xGbB5W�i�ׯ��|2u�02�=�K�3j�o0��p��l��f��[Y_�����\kX�V擴�kͮx�]�����ݮ��������ZS��ge���r�Li����7\�XH:�ܗ��K� ��j A�I���y,�;�sM]����JL�\D	sߓ=�P�#8��8}�
�|�q�-�T�7��$�$PX��JK�3gB`�Z.�f,�R?�-g��<���};6������G����I�����ԑ�K�E���������JLa���"LT��(��t5�B����tg�)pe�L:��U�kn'>� ���L���:�x�l
���LO� ,�'���_:�z�_��8�W� T�<괯��ȝʱ�[�,5��R!��(0�h��q�a�V덾�����l�t><Ho!�|�,���E��0q��2�_&A���p������z��KAK(���Vx�ˇ�����$a��J��_^Ʊ��r�/�Vp��~������{�1���M �N�L�*��iٜ�j�IL���x�����zp�W=����&�2]:�T�BfQr'+0�+��H���O�A2�o���I�tr���ߥ���~�4��掳]�ڮh��<p�`�|yy1�1�N�:C�q?��5s�2��eH�d���ղ�^�7p�_Q,�k�� w���$���܍mݘG�>�ttw��	�ܾ��FR `�5,�[�7�����?n���֠��n�N�~M%K->���#�YN�v�BvFI{h����r���vw_��"܎��#WX��d~)��,-����!d/����W��?�S7�Stc�N��j<���G�S�%��zܞ]���;19y����}����}�
�$S`���e
u[{_�"1��Y��?vQ��v.���D))�]��|e���.Q$V��"w
���Z=��q�eK�x���_iUH��/�~"V�}(⅟�3�o^��>to�9>������������MLl;H��f��G�l��M���RՀvTd�j88�{��5�ҩ&������.��*�.Ê ���>M!߱!w(s:�j�����)��|���D.�9��{��w��EԍHmQ�8��(>�dV0,������Ǖ.�n9�Z�	sh�����f�z��HRZ�_��Uى~yV�L}k&Ο�g��w���2�}�u��W�%y�m���c{���l�����"���|��@@�Q�e>l����:�^�|^���,6�h������K�1��Vݖ��S+�rv���I�ۨp�Ǟ��L]�	��s=|��)z��0G ��BKß�Ά.�ƙ)��Z����ŭ���dn������%�Z��M�W�)K6.�%�t8�5�M�9�����g'GNH�|��y��9���I�.5Ps�J}+B>��]��vfO���F��|�XQ�'�$
�4�����\�Е�dᬕ�zB�#�dK�AyS��"Z�۫�)�0�����0�χ�RZ��u�L'�Y&�J+!w��q�E�*O7rlI&��щ��@���,nA*K�)���0��`�x���.{r X<Rq�������wU���ZvV8����Aa�P�т�ҹ�����@q���)2�� �� s���<�����#��m9���޾����;��p�Oklu��Z+'�4�Z����ڂ�ͽ}綨]�2�z��;����sb�@�ԮG/W�:�әܚ�n�-��Z䆡�������p�)6�]���<Z�O~����<�;w�q�bмk�;ۤ�>ڈ��$]���L�˗���)~A�>�b��ՠ0�F�M߈x��f�;��Q3��"�<�I^�xi��������ؾ��<��,.������f�I�m�=`�)�KmS�C[��3�Y�{�bin>�4��lķ�|\�����0�0ug|>��\��Ϭ��d�jiQ���+�~�B �f+��t�)�-��&��7".�>�ʳ-�)T(͚^�lɲ���)8��v�p��������z��1�=f���Lt?��uLm|{T��Ќ�il�K05�Gfi$n�h)(c���Bܜi#�=}��zV�=�E�m�J<n�*��7������v�9N%�4�|�����4���ʊ*�:V�)��-����)/ґ��#�TV��ǴU�Y� b�X$/��'�ϫ}x�zkvf&�|�DÙ��Fw͌��:n���Y!V��H��8q���X�>H���E"�`���;���� �>5�ף�8�n�&�G�oľ��8�yK,-���F���zt�F<��O���3g� T�-��s�8E:�������7ą�ML5`�P����x�f��]��_��8W��bl�-NG\�(6��x-���Ħ��*�ydCO3>��L�9x)�0���Pl�4�L5R9�����A����L%�%����������+�E?�1�&�b&CX���7��= ��Ҕ��%�BX
*���"坝��N�s2�3�^eH�7'8�!�/Mƻ�>�#�G������#B��H��鹿[0�� ��]B���~;8��eּ�Rvs����/#r�΋$�~�������-q�G��xdr�ֆ+��Sl��֛���.'�ے�DKQrF�-���(7�Z�y�o�����,p���m߫�܏�fץ/��������Ӿ/3��,�g-ꉈ�<W�����ګ�VkW��g8���ҟ[���x��<��_5��>"�
�G�����jq��z��7V80��l�<�@?w��I�[����q�MS 
ܚ�xh]��V�|�?�1�}:ⷿ��kR$J��K��m^�C_���܊|��M�i�.�|�mU���ʐ�3wWBk�&*�i��h����SS�������Է͖ں1\Xn'c��5]%.J)x��;���9���TUVy9�i��+�k�J�<y�V{5�v�Ŷ��%=5����OA���T	��0d>�V�+���Q3��*G�e�"�@�����+[� _�]%��1.am|
~Byƫ�{�˃�V,i��U��ݴ������]�fn�8v����p�O�z<��|�(�}z�}ro�{j_�۳/��\<��g�Ё/�g��l�ܱ'Vfĉ׎���l@ړ@bV!M�C����͘���#�U�������7���;��Bœ�S~����\1�
�&��8׫�M���)[��K�.A�-�-�&(���\-nϖ��հ
n����O���[�˧�)eZX�����c�t=��YB�/���j{�������&�L.�gѩ���`��3#�D����4?��?��x�Qю�����=d���"�����3�����66�P��#U��B�,ȿkk���A71�QT`���3�Z��R�H�дr%@�$]ϴƷm �\�?k:4�;���>MG+ϸ&X���]��;M��;e8��-���㳼wҰ�G�lx�d�1���!L'�:k�U��+?]�ݥ/�o��U�j"�t�9�=GܚN��mҼ��<���&5�"AU#�L�p��:B�S[֊�7mm�3�;cvZYp��0�5c���r+堈Hwv����F��7�d~��,	-C���.�C��٢Qk�����{�C#gS�,�`�-!NPm�w�1�ђ��ȴ�OF-#��X��t��*LCܽ)ϵ厸1��f���sq�c|b&&&o��ܼ��(	\1��)�$t�ɘ�ΛS��G����E�S�f֢�'a2ǈ��|.�-���c;lmY}��4㭇*_g1�kgo��V��c���'�L��SV=��l����r�1�L�R���]��x��N&n�������Áe���ZY�,8B#�_�J��iz©��`��W
�VЦ�eAϖE��"��w>b����6�4�,�*8xS�ƒ�tI&�6A*=���&"����K��V    IEND�B`�PK   l�WW#l��  �     jsons/user_defined.json���n�6�_���Z��D)w�6Nj;A�"(t��B��+Y����R��i�a8���5��~����n��3o�U�W���Q�7������F�`@_�|�{g�?�Yf_�g�m�.f�zP��՗��Ӄ�kq2�x;��RͳXTI�Y�~���ϳ|YȬd1�I�t�q6Ϗ��A���/�z���q^Wu�>�5_�s��Y4U��{��u^��mv7k��=`1�z��ު�~��I*��1������AO�Y��}W�����ھgzQo��T�!a�!������������o��r5���jq{���%>`�*��o%p�	J�  B���e��F_âGxtJ PB�(9 �$N�� E	)� PB�"W�r�K���""����_��q���DB@p�c�MД\[>�)�#�9��LU�n��K.LY�|[���AI8Xnj��H	���)�WF�(���5�Z9��ղ����Qq�e��sܑ�)r~J�9^���ڤ�s���ͻ)�/q�{�'|d��[���ra�VJ_xK�Jc���ȁ��^�������ϗ��|}��)V���d����sl��o*�f��p\*�f�ι9@,_̦GW����	�Ń3��#��M����{������Ե;����fܹmC�_�s��!�����ס�g2k�o�:�#�4�9��P�����%0��J��̑�Kx�#H���#$2d��S�:���c9�,	R��f?1X,?��/�#$���Y,}4��Xz"ſ��� ������$|��s��E�n��0�}�J&+UmU�ϚBM֪��n�R�X�BX�QZ*?i�g����(̀U���ޡ�u�����W�Q��n� 8)H.��$A$�ر`m��w*��M�-[SS� N X���' �5�i�� ���C| _}�֨C����twHN �[Qs�)��|~���12�f6#�9h��X�8���ۇPK
   l�WW5O*@?B  �{                  cirkitFile.jsonPK
   �WWMYMVx�  d�  /             lB  images/010d914f-59de-439a-af91-012b754a10f1.pngPK
   O�WW�.�ɭ � /             13 images/946c31b1-53e3-4800-acb1-710e2b91d3be.pngPK
   <�WW/m�DE! ! /             +@ images/ba63f8f6-a854-4b7a-ba91-7c7ad061d88e.pngPK
   l�WW#l��  �               �a jsons/user_defined.jsonPK      �  �e   